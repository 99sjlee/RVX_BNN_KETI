`default_nettype wire
module BundleBridgeNexus_13(
  output  auto_out
);
  wire  outputs_0 = 1'h0;
  assign auto_out = outputs_0;
endmodule