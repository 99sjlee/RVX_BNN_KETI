// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_126
`define RVX_GDEF_126

`define RVX_GDEF_123 6
`define RVX_GDEF_207 8
`define RVX_GDEF_298 3
`define RVX_GDEF_236 1

`define RVX_GDEF_093 (32'h 0)
`define RVX_GDEF_101 (32'h 8)
`define RVX_GDEF_169 (32'h 10)
`define RVX_GDEF_230 (32'h 18)
`define RVX_GDEF_032 (32'h 20)

`define RVX_GDEF_117 (`RVX_GDEF_093)
`define RVX_GDEF_033 (`RVX_GDEF_101)
`define RVX_GDEF_049 (`RVX_GDEF_169)
`define RVX_GDEF_146 (`RVX_GDEF_230)
`define RVX_GDEF_374 (`RVX_GDEF_032)

`define RVX_GDEF_107 5
`define RVX_GDEF_380 0
`define RVX_GDEF_147 9
`define RVX_GDEF_315 3
`define RVX_GDEF_148 7
`define RVX_GDEF_264 24

`define RVX_GDEF_062 32
`define RVX_GDEF_078 0

`define RVX_GDEF_051 32
`define RVX_GDEF_135 0

`define RVX_GDEF_058 32
`define RVX_GDEF_342 0

`define RVX_GDEF_040 32
`define RVX_GDEF_401 0

`endif