// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_254
`define RVX_GDEF_254

`define RVX_GDEF_234 6
`define RVX_GDEF_133 8
`define RVX_GDEF_188 3
`define RVX_GDEF_375 1

`define RVX_GDEF_177 (32'h 0)
`define RVX_GDEF_201 (32'h 8)
`define RVX_GDEF_249 (32'h 10)
`define RVX_GDEF_141 (32'h 18)
`define RVX_GDEF_042 (32'h 20)
`define RVX_GDEF_299 (32'h 28)

`define RVX_GDEF_109 (`RVX_GDEF_177)
`define RVX_GDEF_258 (`RVX_GDEF_201)
`define RVX_GDEF_312 (`RVX_GDEF_249)
`define RVX_GDEF_079 (`RVX_GDEF_141)
`define RVX_GDEF_417 (`RVX_GDEF_042)
`define RVX_GDEF_371 (`RVX_GDEF_299)

`define RVX_GDEF_284 8
`define RVX_GDEF_358 0
`define RVX_GDEF_038 1
`define RVX_GDEF_433 2
`define RVX_GDEF_198 4
`define RVX_GDEF_430 8
`define RVX_GDEF_212 16
`define RVX_GDEF_296 32
`define RVX_GDEF_192 64
`define RVX_GDEF_225 128
`define RVX_GDEF_422 0
`define RVX_GDEF_167 1
`define RVX_GDEF_246 2
`define RVX_GDEF_335 3
`define RVX_GDEF_337 4
`define RVX_GDEF_149 5
`define RVX_GDEF_172 6
`define RVX_GDEF_130 7
`define RVX_GDEF_137 0

`define RVX_GDEF_037 5
`define RVX_GDEF_046 0
`define RVX_GDEF_215 1
`define RVX_GDEF_039 2
`define RVX_GDEF_285 4
`define RVX_GDEF_309 8
`define RVX_GDEF_400 16
`define RVX_GDEF_199 0
`define RVX_GDEF_410 1
`define RVX_GDEF_307 2
`define RVX_GDEF_151 3
`define RVX_GDEF_083 4
`define RVX_GDEF_229 0

`define RVX_GDEF_061 8
`define RVX_GDEF_187 0

`define RVX_GDEF_368 32
`define RVX_GDEF_182 0

`define RVX_GDEF_399 32
`define RVX_GDEF_302 0

`define RVX_GDEF_291 7
`define RVX_GDEF_317 0

`endif