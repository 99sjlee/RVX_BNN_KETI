// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_253
`define RVX_GDEF_253

`define RVX_GDEF_294 6
`define RVX_GDEF_115 8
`define RVX_GDEF_025 3
`define RVX_GDEF_419 1

`define RVX_GDEF_170 (32'h 0)
`define RVX_GDEF_322 (32'h 8)
`define RVX_GDEF_206 (32'h 10)
`define RVX_GDEF_204 (32'h 18)
`define RVX_GDEF_349 (32'h 20)

`define RVX_GDEF_168 (`RVX_GDEF_170)
`define RVX_GDEF_134 (`RVX_GDEF_322)
`define RVX_GDEF_289 (`RVX_GDEF_206)
`define RVX_GDEF_373 (`RVX_GDEF_204)
`define RVX_GDEF_183 (`RVX_GDEF_349)

`define RVX_GDEF_184 1
`define RVX_GDEF_310 0
`define RVX_GDEF_277 1
`define RVX_GDEF_343 0
`define RVX_GDEF_431 0

`define RVX_GDEF_075 32
`define RVX_GDEF_159 0

`define RVX_GDEF_222 32
`define RVX_GDEF_108 0

`define RVX_GDEF_153 32
`define RVX_GDEF_043 0

`define RVX_GDEF_233 32
`define RVX_GDEF_268 0

`define RVX_GDEF_248 32
`define RVX_GDEF_171 0

`endif