`default_nettype wire
module OptimizationBarrier_42(
  input  [2:0] io_x,
  output [2:0] io_y
);
  assign io_y = io_x;
endmodule