`default_nettype wire
module CSRFile(
  input         clock,
  input         reset,
  input         io_ungated_clock,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  input         io_hartid,
  input  [11:0] io_rw_addr,
  input  [2:0]  io_rw_cmd,
  output [31:0] io_rw_rdata,
  input  [31:0] io_rw_wdata,
  input  [31:0] io_decode_0_inst,
  output        io_decode_0_fp_illegal,
  output        io_decode_0_fp_csr,
  output        io_decode_0_rocc_illegal,
  output        io_decode_0_read_illegal,
  output        io_decode_0_write_illegal,
  output        io_decode_0_write_flush,
  output        io_decode_0_system_illegal,
  output        io_csr_stall,
  output        io_eret,
  output        io_singleStep,
  output        io_status_debug,
  output        io_status_cease,
  output        io_status_wfi,
  output [31:0] io_status_isa,
  output [1:0]  io_status_dprv,
  output        io_status_dv,
  output [1:0]  io_status_prv,
  output        io_status_v,
  output        io_status_sd,
  output [22:0] io_status_zero2,
  output        io_status_mpv,
  output        io_status_gva,
  output        io_status_mbe,
  output        io_status_sbe,
  output [1:0]  io_status_sxl,
  output [1:0]  io_status_uxl,
  output        io_status_sd_rv32,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_vs,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_ube,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output        io_ptbr_mode,
  output [21:0] io_ptbr_ppn,
  output [31:0] io_evec,
  input         io_exception,
  input         io_retire,
  input  [31:0] io_cause,
  input  [31:0] io_pc,
  input  [31:0] io_tval,
  input         io_gva,
  output [31:0] io_time,
  output [2:0]  io_fcsr_rm,
  input         io_fcsr_flags_valid,
  input  [4:0]  io_fcsr_flags_bits,
  output        io_interrupt,
  output [31:0] io_interrupt_cause,
  output        io_bp_0_control_action,
  output [1:0]  io_bp_0_control_tmatch,
  output        io_bp_0_control_m,
  output        io_bp_0_control_s,
  output        io_bp_0_control_u,
  output        io_bp_0_control_x,
  output        io_bp_0_control_w,
  output        io_bp_0_control_r,
  output [31:0] io_bp_0_address,
  output        io_pmp_0_cfg_l,
  output [1:0]  io_pmp_0_cfg_a,
  output        io_pmp_0_cfg_x,
  output        io_pmp_0_cfg_w,
  output        io_pmp_0_cfg_r,
  output [29:0] io_pmp_0_addr,
  output [31:0] io_pmp_0_mask,
  output        io_pmp_1_cfg_l,
  output [1:0]  io_pmp_1_cfg_a,
  output        io_pmp_1_cfg_x,
  output        io_pmp_1_cfg_w,
  output        io_pmp_1_cfg_r,
  output [29:0] io_pmp_1_addr,
  output [31:0] io_pmp_1_mask,
  output        io_pmp_2_cfg_l,
  output [1:0]  io_pmp_2_cfg_a,
  output        io_pmp_2_cfg_x,
  output        io_pmp_2_cfg_w,
  output        io_pmp_2_cfg_r,
  output [29:0] io_pmp_2_addr,
  output [31:0] io_pmp_2_mask,
  output        io_pmp_3_cfg_l,
  output [1:0]  io_pmp_3_cfg_a,
  output        io_pmp_3_cfg_x,
  output        io_pmp_3_cfg_w,
  output        io_pmp_3_cfg_r,
  output [29:0] io_pmp_3_addr,
  output [31:0] io_pmp_3_mask,
  output        io_pmp_4_cfg_l,
  output [1:0]  io_pmp_4_cfg_a,
  output        io_pmp_4_cfg_x,
  output        io_pmp_4_cfg_w,
  output        io_pmp_4_cfg_r,
  output [29:0] io_pmp_4_addr,
  output [31:0] io_pmp_4_mask,
  output        io_pmp_5_cfg_l,
  output [1:0]  io_pmp_5_cfg_a,
  output        io_pmp_5_cfg_x,
  output        io_pmp_5_cfg_w,
  output        io_pmp_5_cfg_r,
  output [29:0] io_pmp_5_addr,
  output [31:0] io_pmp_5_mask,
  output        io_pmp_6_cfg_l,
  output [1:0]  io_pmp_6_cfg_a,
  output        io_pmp_6_cfg_x,
  output        io_pmp_6_cfg_w,
  output        io_pmp_6_cfg_r,
  output [29:0] io_pmp_6_addr,
  output [31:0] io_pmp_6_mask,
  output        io_pmp_7_cfg_l,
  output [1:0]  io_pmp_7_cfg_a,
  output        io_pmp_7_cfg_x,
  output        io_pmp_7_cfg_w,
  output        io_pmp_7_cfg_r,
  output [29:0] io_pmp_7_addr,
  output [31:0] io_pmp_7_mask,
  output        io_inhibit_cycle,
  input  [31:0] io_inst_0,
  output        io_trace_0_valid,
  output [31:0] io_trace_0_iaddr,
  output [31:0] io_trace_0_insn,
  output        io_trace_0_exception,
  output [31:0] io_customCSRs_0_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] reg_mstatus_prv;
  reg  reg_mstatus_gva;
  reg  reg_mstatus_tsr;
  reg  reg_mstatus_tw;
  reg  reg_mstatus_tvm;
  reg  reg_mstatus_mxr;
  reg  reg_mstatus_sum;
  reg  reg_mstatus_mprv;
  reg [1:0] reg_mstatus_fs;
  reg [1:0] reg_mstatus_mpp;
  reg  reg_mstatus_spp;
  reg  reg_mstatus_mpie;
  reg  reg_mstatus_spie;
  reg  reg_mstatus_mie;
  reg  reg_mstatus_sie;
  wire  system_insn = io_rw_cmd == 3'h4;
  wire [31:0] _T_330 = {io_rw_addr, 20'h0};
  wire [31:0] decoded_plaInput = 32'h73 | _T_330;
  wire [31:0] decoded_invInputs = ~decoded_plaInput;
  wire  decoded_andMatrixInput_0 = decoded_invInputs[20];
  wire  decoded_andMatrixInput_1 = decoded_invInputs[21];
  wire  decoded_andMatrixInput_2 = decoded_invInputs[22];
  wire  decoded_andMatrixInput_3 = decoded_invInputs[23];
  wire  decoded_andMatrixInput_4 = decoded_invInputs[24];
  wire  decoded_andMatrixInput_5 = decoded_invInputs[25];
  wire  decoded_andMatrixInput_6 = decoded_invInputs[26];
  wire  decoded_andMatrixInput_7 = decoded_invInputs[27];
  wire  decoded_andMatrixInput_8 = decoded_invInputs[28];
  wire  decoded_andMatrixInput_9 = decoded_invInputs[29];
  wire  decoded_andMatrixInput_10 = decoded_invInputs[30];
  wire  decoded_andMatrixInput_11 = decoded_invInputs[31];
  wire [5:0] decoded_lo = {decoded_andMatrixInput_6,decoded_andMatrixInput_7,decoded_andMatrixInput_8,
    decoded_andMatrixInput_9,decoded_andMatrixInput_10,decoded_andMatrixInput_11};
  wire [11:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4,decoded_andMatrixInput_5,decoded_lo};
  wire  _decoded_T_1 = &_decoded_T;
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_T_1;
  wire  decoded_andMatrixInput_0_1 = decoded_plaInput[20];
  wire [11:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4,decoded_andMatrixInput_5,decoded_lo};
  wire  _decoded_T_3 = &_decoded_T_2;
  wire  _decoded_orMatrixOutputs_T_5 = |_decoded_T_3;
  wire  decoded_andMatrixInput_0_2 = decoded_plaInput[0];
  wire  decoded_andMatrixInput_7_2 = decoded_plaInput[28];
  wire [9:0] _decoded_T_4 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_2,decoded_andMatrixInput_3,
    decoded_andMatrixInput_4,decoded_andMatrixInput_5,decoded_andMatrixInput_6,decoded_andMatrixInput_7,
    decoded_andMatrixInput_7_2,decoded_andMatrixInput_10,decoded_andMatrixInput_11};
  wire  _decoded_T_5 = &_decoded_T_4;
  wire  decoded_andMatrixInput_0_6 = decoded_plaInput[30];
  wire [1:0] _decoded_T_12 = {decoded_andMatrixInput_0_6,decoded_andMatrixInput_11};
  wire  _decoded_T_13 = &_decoded_T_12;
  wire [1:0] _decoded_orMatrixOutputs_T_3 = {_decoded_T_5,_decoded_T_13};
  wire  _decoded_orMatrixOutputs_T_4 = |_decoded_orMatrixOutputs_T_3;
  wire  decoded_andMatrixInput_0_5 = decoded_plaInput[22];
  wire  decoded_andMatrixInput_7_5 = decoded_plaInput[29];
  wire [9:0] _decoded_T_10 = {decoded_andMatrixInput_0_5,decoded_andMatrixInput_3,decoded_andMatrixInput_4,
    decoded_andMatrixInput_5,decoded_andMatrixInput_6,decoded_andMatrixInput_7,decoded_andMatrixInput_7_2,
    decoded_andMatrixInput_7_5,decoded_andMatrixInput_10,decoded_andMatrixInput_11};
  wire  _decoded_T_11 = &_decoded_T_10;
  wire  _decoded_orMatrixOutputs_T_2 = |_decoded_T_11;
  wire [9:0] _decoded_T_6 = {decoded_andMatrixInput_0_5,decoded_andMatrixInput_3,decoded_andMatrixInput_4,
    decoded_andMatrixInput_5,decoded_andMatrixInput_6,decoded_andMatrixInput_7,decoded_andMatrixInput_7_2,
    decoded_andMatrixInput_9,decoded_andMatrixInput_10,decoded_andMatrixInput_11};
  wire  _decoded_T_7 = &_decoded_T_6;
  wire  _decoded_orMatrixOutputs_T_1 = |_decoded_T_7;
  wire  decoded_andMatrixInput_1_4 = decoded_plaInput[1];
  wire  decoded_andMatrixInput_2_4 = decoded_invInputs[2];
  wire  decoded_andMatrixInput_3_4 = decoded_invInputs[3];
  wire  decoded_andMatrixInput_4_4 = decoded_plaInput[4];
  wire  decoded_andMatrixInput_5_4 = decoded_plaInput[5];
  wire  decoded_andMatrixInput_6_4 = decoded_plaInput[6];
  wire  decoded_andMatrixInput_7_4 = decoded_invInputs[7];
  wire  decoded_andMatrixInput_8_4 = decoded_invInputs[8];
  wire  decoded_andMatrixInput_9_4 = decoded_invInputs[9];
  wire  decoded_andMatrixInput_10_2 = decoded_plaInput[25];
  wire [7:0] decoded_lo_4 = {decoded_andMatrixInput_9_4,decoded_andMatrixInput_10_2,decoded_andMatrixInput_6,
    decoded_andMatrixInput_7,decoded_andMatrixInput_7_2,decoded_andMatrixInput_9,decoded_andMatrixInput_10,
    decoded_andMatrixInput_11};
  wire [16:0] _decoded_T_8 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_1_4,decoded_andMatrixInput_2_4,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_4,decoded_andMatrixInput_5_4,decoded_andMatrixInput_6_4,
    decoded_andMatrixInput_7_4,decoded_andMatrixInput_8_4,decoded_lo_4};
  wire  _decoded_T_9 = &_decoded_T_8;
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_9;
  wire [8:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_5,
    _decoded_orMatrixOutputs_T_4,_decoded_orMatrixOutputs_T_2,_decoded_orMatrixOutputs_T_1,_decoded_orMatrixOutputs_T,1'h0
    ,2'h0};
  wire [8:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[8],decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6
    ],decoded_orMatrixOutputs[5],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],
    decoded_orMatrixOutputs[1],decoded_orMatrixOutputs[0]};
  wire  insn_ret = system_insn & decoded_invMatrixOutputs[6];
  reg [1:0] reg_dcsr_prv;
  wire [1:0] _GEN_236 = io_rw_addr[10] & io_rw_addr[7] ? reg_dcsr_prv : reg_mstatus_mpp;
  wire [1:0] ret_prv = ~io_rw_addr[9] ? {{1'd0}, reg_mstatus_spp} : _GEN_236;
  wire  insn_call = system_insn & decoded_invMatrixOutputs[8];
  wire  insn_break = system_insn & decoded_invMatrixOutputs[7];
  wire  _exception_T = insn_call | insn_break;
  wire  exception = insn_call | insn_break | io_exception;
  reg  reg_singleStepped;
  wire [3:0] _GEN_34 = {{2'd0}, reg_mstatus_prv};
  wire [3:0] _cause_T_4 = 4'h8 + _GEN_34;
  wire [31:0] _cause_T_5 = insn_break ? 32'h3 : io_cause;
  wire [31:0] cause = insn_call ? {{28'd0}, _cause_T_4} : _cause_T_5;
  wire [7:0] cause_lsbs = cause[7:0];
  wire  _causeIsDebugInt_T_1 = cause_lsbs == 8'he;
  wire  causeIsDebugInt = cause[31] & cause_lsbs == 8'he;
  wire  _causeIsDebugTrigger_T_1 = ~cause[31];
  wire  causeIsDebugTrigger = ~cause[31] & _causeIsDebugInt_T_1;
  reg  reg_dcsr_ebreakm;
  reg  reg_dcsr_ebreaks;
  reg  reg_dcsr_ebreaku;
  wire [3:0] _causeIsDebugBreak_T_3 = {reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  wire [3:0] _causeIsDebugBreak_T_4 = _causeIsDebugBreak_T_3 >> reg_mstatus_prv;
  wire  causeIsDebugBreak = _causeIsDebugTrigger_T_1 & insn_break & _causeIsDebugBreak_T_4[0];
  reg  reg_debug;
  wire  trapToDebug = reg_singleStepped | causeIsDebugInt | causeIsDebugTrigger | causeIsDebugBreak | reg_debug;
  wire  _T_397 = ~reg_debug;
  wire [1:0] _GEN_56 = ~reg_debug ? 2'h3 : reg_mstatus_prv;
  wire  _delegate_T = reg_mstatus_prv <= 2'h1;
  reg [31:0] reg_mideleg;
  wire [31:0] read_mideleg = reg_mideleg & 32'h222;
  wire [31:0] _delegate_T_3 = read_mideleg >> cause_lsbs;
  reg [31:0] reg_medeleg;
  wire [31:0] read_medeleg = reg_medeleg & 32'hf0b55d;
  wire [31:0] _delegate_T_5 = read_medeleg >> cause_lsbs;
  wire  _delegate_T_7 = cause[31] ? _delegate_T_3[0] : _delegate_T_5[0];
  wire  delegate = reg_mstatus_prv <= 2'h1 & _delegate_T_7;
  wire [1:0] _GEN_75 = delegate ? 2'h1 : 2'h3;
  wire [1:0] _GEN_150 = trapToDebug ? _GEN_56 : _GEN_75;
  wire [1:0] _GEN_187 = exception ? _GEN_150 : reg_mstatus_prv;
  wire [1:0] new_prv = insn_ret ? ret_prv : _GEN_187;
  reg [2:0] reg_dcsr_cause;
  reg  reg_dcsr_step;
  reg [31:0] reg_dpc;
  reg [31:0] reg_dscratch0;
  reg  reg_bp_0_control_dmode;
  reg  reg_bp_0_control_action;
  reg [1:0] reg_bp_0_control_tmatch;
  reg  reg_bp_0_control_m;
  reg  reg_bp_0_control_s;
  reg  reg_bp_0_control_u;
  reg  reg_bp_0_control_x;
  reg  reg_bp_0_control_w;
  reg  reg_bp_0_control_r;
  reg [31:0] reg_bp_0_address;
  reg  reg_pmp_0_cfg_l;
  reg [1:0] reg_pmp_0_cfg_a;
  reg  reg_pmp_0_cfg_x;
  reg  reg_pmp_0_cfg_w;
  reg  reg_pmp_0_cfg_r;
  reg [29:0] reg_pmp_0_addr;
  reg  reg_pmp_1_cfg_l;
  reg [1:0] reg_pmp_1_cfg_a;
  reg  reg_pmp_1_cfg_x;
  reg  reg_pmp_1_cfg_w;
  reg  reg_pmp_1_cfg_r;
  reg [29:0] reg_pmp_1_addr;
  reg  reg_pmp_2_cfg_l;
  reg [1:0] reg_pmp_2_cfg_a;
  reg  reg_pmp_2_cfg_x;
  reg  reg_pmp_2_cfg_w;
  reg  reg_pmp_2_cfg_r;
  reg [29:0] reg_pmp_2_addr;
  reg  reg_pmp_3_cfg_l;
  reg [1:0] reg_pmp_3_cfg_a;
  reg  reg_pmp_3_cfg_x;
  reg  reg_pmp_3_cfg_w;
  reg  reg_pmp_3_cfg_r;
  reg [29:0] reg_pmp_3_addr;
  reg  reg_pmp_4_cfg_l;
  reg [1:0] reg_pmp_4_cfg_a;
  reg  reg_pmp_4_cfg_x;
  reg  reg_pmp_4_cfg_w;
  reg  reg_pmp_4_cfg_r;
  reg [29:0] reg_pmp_4_addr;
  reg  reg_pmp_5_cfg_l;
  reg [1:0] reg_pmp_5_cfg_a;
  reg  reg_pmp_5_cfg_x;
  reg  reg_pmp_5_cfg_w;
  reg  reg_pmp_5_cfg_r;
  reg [29:0] reg_pmp_5_addr;
  reg  reg_pmp_6_cfg_l;
  reg [1:0] reg_pmp_6_cfg_a;
  reg  reg_pmp_6_cfg_x;
  reg  reg_pmp_6_cfg_w;
  reg  reg_pmp_6_cfg_r;
  reg [29:0] reg_pmp_6_addr;
  reg  reg_pmp_7_cfg_l;
  reg [1:0] reg_pmp_7_cfg_a;
  reg  reg_pmp_7_cfg_x;
  reg  reg_pmp_7_cfg_w;
  reg  reg_pmp_7_cfg_r;
  reg [29:0] reg_pmp_7_addr;
  reg [31:0] reg_mie;
  reg  reg_mip_seip;
  reg  reg_mip_stip;
  reg  reg_mip_ssip;
  reg [31:0] reg_mepc;
  reg [31:0] reg_mcause;
  reg [31:0] reg_mtval;
  reg [31:0] reg_mscratch;
  reg [31:0] reg_mtvec;
  reg [31:0] reg_mcounteren;
  wire [31:0] read_mcounteren = reg_mcounteren & 32'h7;
  reg [31:0] reg_scounteren;
  wire [31:0] read_scounteren = reg_scounteren & 32'h7;
  wire [15:0] _read_hvip_T = {4'h0,2'h0,reg_mip_seip,1'h0,2'h0,reg_mip_stip,1'h0,2'h0,reg_mip_ssip,1'h0};
  reg [31:0] reg_sepc;
  reg [31:0] reg_scause;
  reg [31:0] reg_stval;
  reg [31:0] reg_sscratch;
  reg [31:0] reg_stvec;
  reg  reg_satp_mode;
  reg [21:0] reg_satp_ppn;
  reg  reg_wfi;
  reg [4:0] reg_fflags;
  reg [2:0] reg_frm;
  reg [2:0] reg_mcountinhibit;
  wire  x79 = reg_mcountinhibit[2];
  reg [5:0] small_;
  wire [5:0] _GEN_35 = {{5'd0}, io_retire};
  wire [6:0] nextSmall = small_ + _GEN_35;
  wire  _T_14 = ~x79;
  wire [6:0] _GEN_0 = ~x79 ? nextSmall : {{1'd0}, small_};
  reg [57:0] large_;
  wire [57:0] _large_r_T_1 = large_ + 58'h1;
  wire [57:0] _GEN_1 = nextSmall[6] & _T_14 ? _large_r_T_1 : large_;
  wire [63:0] value = {large_,small_};
  wire  x86 = ~io_csr_stall;
  reg [5:0] small_1;
  wire [5:0] _GEN_40 = {{5'd0}, x86};
  wire [6:0] nextSmall_1 = small_1 + _GEN_40;
  wire  _T_15 = ~reg_mcountinhibit[0];
  wire [6:0] _GEN_2 = ~reg_mcountinhibit[0] ? nextSmall_1 : {{1'd0}, small_1};
  reg [57:0] large_1;
  wire [57:0] _large_r_T_3 = large_1 + 58'h1;
  wire [57:0] _GEN_3 = nextSmall_1[6] & _T_15 ? _large_r_T_3 : large_1;
  wire [63:0] value_1 = {large_1,small_1};
  wire  mip_seip = reg_mip_seip | io_interrupts_seip;
  wire [7:0] read_mip_lo = {io_interrupts_mtip,1'h0,reg_mip_stip,1'h0,io_interrupts_msip,1'h0,reg_mip_ssip,1'h0};
  wire [15:0] _read_mip_T = {4'h0,io_interrupts_meip,1'h0,mip_seip,1'h0,read_mip_lo};
  wire [15:0] read_mip = _read_mip_T & 16'haaa;
  wire [31:0] _GEN_41 = {{16'd0}, read_mip};
  wire [31:0] pending_interrupts = _GEN_41 & reg_mie;
  wire [14:0] d_interrupts = {io_interrupts_debug, 14'h0};
  wire [31:0] _m_interrupts_T_3 = ~pending_interrupts;
  wire [31:0] _m_interrupts_T_4 = _m_interrupts_T_3 | read_mideleg;
  wire [31:0] _m_interrupts_T_5 = ~_m_interrupts_T_4;
  wire [31:0] m_interrupts = _delegate_T | reg_mstatus_mie ? _m_interrupts_T_5 : 32'h0;
  wire [31:0] _s_interrupts_T_6 = pending_interrupts & read_mideleg;
  wire [31:0] s_interrupts = reg_mstatus_prv < 2'h1 | reg_mstatus_prv == 2'h1 & reg_mstatus_sie ? _s_interrupts_T_6 : 32'h0
    ;
  wire  _any_T_78 = d_interrupts[14] | d_interrupts[13] | d_interrupts[12] | d_interrupts[11] | d_interrupts[3] |
    d_interrupts[7] | d_interrupts[9] | d_interrupts[1] | d_interrupts[5] | d_interrupts[10] | d_interrupts[2] |
    d_interrupts[6] | d_interrupts[8] | d_interrupts[0] | d_interrupts[4] | m_interrupts[15];
  wire  _any_T_93 = _any_T_78 | m_interrupts[14] | m_interrupts[13] | m_interrupts[12] | m_interrupts[11] | m_interrupts
    [3] | m_interrupts[7] | m_interrupts[9] | m_interrupts[1] | m_interrupts[5] | m_interrupts[10] | m_interrupts[2] |
    m_interrupts[6] | m_interrupts[8] | m_interrupts[0] | m_interrupts[4];
  wire  _any_T_108 = _any_T_93 | s_interrupts[15] | s_interrupts[14] | s_interrupts[13] | s_interrupts[12] |
    s_interrupts[11] | s_interrupts[3] | s_interrupts[7] | s_interrupts[9] | s_interrupts[1] | s_interrupts[5] |
    s_interrupts[10] | s_interrupts[2] | s_interrupts[6] | s_interrupts[8] | s_interrupts[0];
  wire  anyInterrupt = _any_T_108 | s_interrupts[4];
  wire [3:0] _which_T_79 = s_interrupts[0] ? 4'h0 : 4'h4;
  wire [3:0] _which_T_80 = s_interrupts[8] ? 4'h8 : _which_T_79;
  wire [3:0] _which_T_81 = s_interrupts[6] ? 4'h6 : _which_T_80;
  wire [3:0] _which_T_82 = s_interrupts[2] ? 4'h2 : _which_T_81;
  wire [3:0] _which_T_83 = s_interrupts[10] ? 4'ha : _which_T_82;
  wire [3:0] _which_T_84 = s_interrupts[5] ? 4'h5 : _which_T_83;
  wire [3:0] _which_T_85 = s_interrupts[1] ? 4'h1 : _which_T_84;
  wire [3:0] _which_T_86 = s_interrupts[9] ? 4'h9 : _which_T_85;
  wire [3:0] _which_T_87 = s_interrupts[7] ? 4'h7 : _which_T_86;
  wire [3:0] _which_T_88 = s_interrupts[3] ? 4'h3 : _which_T_87;
  wire [3:0] _which_T_89 = s_interrupts[11] ? 4'hb : _which_T_88;
  wire [3:0] _which_T_90 = s_interrupts[12] ? 4'hc : _which_T_89;
  wire [3:0] _which_T_91 = s_interrupts[13] ? 4'hd : _which_T_90;
  wire [3:0] _which_T_92 = s_interrupts[14] ? 4'he : _which_T_91;
  wire [3:0] _which_T_93 = s_interrupts[15] ? 4'hf : _which_T_92;
  wire [3:0] _which_T_94 = m_interrupts[4] ? 4'h4 : _which_T_93;
  wire [3:0] _which_T_95 = m_interrupts[0] ? 4'h0 : _which_T_94;
  wire [3:0] _which_T_96 = m_interrupts[8] ? 4'h8 : _which_T_95;
  wire [3:0] _which_T_97 = m_interrupts[6] ? 4'h6 : _which_T_96;
  wire [3:0] _which_T_98 = m_interrupts[2] ? 4'h2 : _which_T_97;
  wire [3:0] _which_T_99 = m_interrupts[10] ? 4'ha : _which_T_98;
  wire [3:0] _which_T_100 = m_interrupts[5] ? 4'h5 : _which_T_99;
  wire [3:0] _which_T_101 = m_interrupts[1] ? 4'h1 : _which_T_100;
  wire [3:0] _which_T_102 = m_interrupts[9] ? 4'h9 : _which_T_101;
  wire [3:0] _which_T_103 = m_interrupts[7] ? 4'h7 : _which_T_102;
  wire [3:0] _which_T_104 = m_interrupts[3] ? 4'h3 : _which_T_103;
  wire [3:0] _which_T_105 = m_interrupts[11] ? 4'hb : _which_T_104;
  wire [3:0] _which_T_106 = m_interrupts[12] ? 4'hc : _which_T_105;
  wire [3:0] _which_T_107 = m_interrupts[13] ? 4'hd : _which_T_106;
  wire [3:0] _which_T_108 = m_interrupts[14] ? 4'he : _which_T_107;
  wire [3:0] _which_T_109 = m_interrupts[15] ? 4'hf : _which_T_108;
  wire [3:0] _which_T_111 = d_interrupts[4] ? 4'h4 : _which_T_109;
  wire [3:0] _which_T_112 = d_interrupts[0] ? 4'h0 : _which_T_111;
  wire [3:0] _which_T_113 = d_interrupts[8] ? 4'h8 : _which_T_112;
  wire [3:0] _which_T_114 = d_interrupts[6] ? 4'h6 : _which_T_113;
  wire [3:0] _which_T_115 = d_interrupts[2] ? 4'h2 : _which_T_114;
  wire [3:0] _which_T_116 = d_interrupts[10] ? 4'ha : _which_T_115;
  wire [3:0] _which_T_117 = d_interrupts[5] ? 4'h5 : _which_T_116;
  wire [3:0] _which_T_118 = d_interrupts[1] ? 4'h1 : _which_T_117;
  wire [3:0] _which_T_119 = d_interrupts[9] ? 4'h9 : _which_T_118;
  wire [3:0] _which_T_120 = d_interrupts[7] ? 4'h7 : _which_T_119;
  wire [3:0] _which_T_121 = d_interrupts[3] ? 4'h3 : _which_T_120;
  wire [3:0] _which_T_122 = d_interrupts[11] ? 4'hb : _which_T_121;
  wire [3:0] _which_T_123 = d_interrupts[12] ? 4'hc : _which_T_122;
  wire [3:0] _which_T_124 = d_interrupts[13] ? 4'hd : _which_T_123;
  wire [3:0] whichInterrupt = d_interrupts[14] ? 4'he : _which_T_124;
  wire [31:0] _GEN_663 = {{28'd0}, whichInterrupt};
  wire  _io_interrupt_T = ~io_singleStep;
  wire [30:0] pmp_mask_base = {reg_pmp_0_addr,reg_pmp_0_cfg_a[0]};
  wire [30:0] _pmp_mask_T_1 = pmp_mask_base + 31'h1;
  wire [30:0] _pmp_mask_T_2 = ~_pmp_mask_T_1;
  wire [30:0] _pmp_mask_T_3 = pmp_mask_base & _pmp_mask_T_2;
  wire [32:0] _pmp_mask_T_4 = {_pmp_mask_T_3,2'h3};
  wire [30:0] pmp_mask_base_1 = {reg_pmp_1_addr,reg_pmp_1_cfg_a[0]};
  wire [30:0] _pmp_mask_T_6 = pmp_mask_base_1 + 31'h1;
  wire [30:0] _pmp_mask_T_7 = ~_pmp_mask_T_6;
  wire [30:0] _pmp_mask_T_8 = pmp_mask_base_1 & _pmp_mask_T_7;
  wire [32:0] _pmp_mask_T_9 = {_pmp_mask_T_8,2'h3};
  wire [30:0] pmp_mask_base_2 = {reg_pmp_2_addr,reg_pmp_2_cfg_a[0]};
  wire [30:0] _pmp_mask_T_11 = pmp_mask_base_2 + 31'h1;
  wire [30:0] _pmp_mask_T_12 = ~_pmp_mask_T_11;
  wire [30:0] _pmp_mask_T_13 = pmp_mask_base_2 & _pmp_mask_T_12;
  wire [32:0] _pmp_mask_T_14 = {_pmp_mask_T_13,2'h3};
  wire [30:0] pmp_mask_base_3 = {reg_pmp_3_addr,reg_pmp_3_cfg_a[0]};
  wire [30:0] _pmp_mask_T_16 = pmp_mask_base_3 + 31'h1;
  wire [30:0] _pmp_mask_T_17 = ~_pmp_mask_T_16;
  wire [30:0] _pmp_mask_T_18 = pmp_mask_base_3 & _pmp_mask_T_17;
  wire [32:0] _pmp_mask_T_19 = {_pmp_mask_T_18,2'h3};
  wire [30:0] pmp_mask_base_4 = {reg_pmp_4_addr,reg_pmp_4_cfg_a[0]};
  wire [30:0] _pmp_mask_T_21 = pmp_mask_base_4 + 31'h1;
  wire [30:0] _pmp_mask_T_22 = ~_pmp_mask_T_21;
  wire [30:0] _pmp_mask_T_23 = pmp_mask_base_4 & _pmp_mask_T_22;
  wire [32:0] _pmp_mask_T_24 = {_pmp_mask_T_23,2'h3};
  wire [30:0] pmp_mask_base_5 = {reg_pmp_5_addr,reg_pmp_5_cfg_a[0]};
  wire [30:0] _pmp_mask_T_26 = pmp_mask_base_5 + 31'h1;
  wire [30:0] _pmp_mask_T_27 = ~_pmp_mask_T_26;
  wire [30:0] _pmp_mask_T_28 = pmp_mask_base_5 & _pmp_mask_T_27;
  wire [32:0] _pmp_mask_T_29 = {_pmp_mask_T_28,2'h3};
  wire [30:0] pmp_mask_base_6 = {reg_pmp_6_addr,reg_pmp_6_cfg_a[0]};
  wire [30:0] _pmp_mask_T_31 = pmp_mask_base_6 + 31'h1;
  wire [30:0] _pmp_mask_T_32 = ~_pmp_mask_T_31;
  wire [30:0] _pmp_mask_T_33 = pmp_mask_base_6 & _pmp_mask_T_32;
  wire [32:0] _pmp_mask_T_34 = {_pmp_mask_T_33,2'h3};
  wire [30:0] pmp_mask_base_7 = {reg_pmp_7_addr,reg_pmp_7_cfg_a[0]};
  wire [30:0] _pmp_mask_T_36 = pmp_mask_base_7 + 31'h1;
  wire [30:0] _pmp_mask_T_37 = ~_pmp_mask_T_36;
  wire [30:0] _pmp_mask_T_38 = pmp_mask_base_7 & _pmp_mask_T_37;
  wire [32:0] _pmp_mask_T_39 = {_pmp_mask_T_38,2'h3};
  reg [31:0] reg_misa;
  wire [8:0] read_mstatus_lo_lo = {io_status_spp,io_status_mpie,io_status_ube,io_status_spie,io_status_upie,
    io_status_mie,io_status_hie,io_status_sie,io_status_uie};
  wire [21:0] read_mstatus_lo = {io_status_tw,io_status_tvm,io_status_mxr,io_status_sum,io_status_mprv,io_status_xs,
    io_status_fs,io_status_mpp,io_status_vs,read_mstatus_lo_lo};
  wire [64:0] read_mstatus_hi_hi = {io_status_debug,io_status_cease,io_status_wfi,io_status_isa,io_status_dprv,
    io_status_dv,io_status_prv,io_status_v,io_status_sd,io_status_zero2};
  wire [82:0] read_mstatus_hi = {read_mstatus_hi_hi,io_status_mpv,io_status_gva,io_status_mbe,io_status_sbe,
    io_status_sxl,io_status_uxl,io_status_sd_rv32,io_status_zero1,io_status_tsr};
  wire [104:0] _read_mstatus_T = {read_mstatus_hi,read_mstatus_lo};
  wire [31:0] read_mstatus = _read_mstatus_T[31:0];
  wire [6:0] _read_mtvec_T_1 = reg_mtvec[0] ? 7'h7e : 7'h2;
  wire [31:0] _read_mtvec_T_3 = {{25'd0}, _read_mtvec_T_1};
  wire [31:0] _read_mtvec_T_4 = ~_read_mtvec_T_3;
  wire [31:0] read_mtvec = reg_mtvec & _read_mtvec_T_4;
  wire [6:0] _read_stvec_T_1 = reg_stvec[0] ? 7'h7e : 7'h2;
  wire [31:0] _read_stvec_T_3 = {{25'd0}, _read_stvec_T_1};
  wire [31:0] _read_stvec_T_4 = ~_read_stvec_T_3;
  wire [31:0] read_stvec = reg_stvec & _read_stvec_T_4;
  wire [6:0] lo_4 = {reg_bp_0_control_m,1'h0,reg_bp_0_control_s,reg_bp_0_control_u,reg_bp_0_control_x,reg_bp_0_control_w
    ,reg_bp_0_control_r};
  wire [31:0] _T_16 = {4'h2,reg_bp_0_control_dmode,14'h400,reg_bp_0_control_action,1'h0,2'h0,reg_bp_0_control_tmatch,
    lo_4};
  wire [31:0] _T_18 = ~reg_mepc;
  wire [1:0] _T_20 = reg_misa[2] ? 2'h1 : 2'h3;
  wire [31:0] _GEN_664 = {{30'd0}, _T_20};
  wire [31:0] _T_21 = _T_18 | _GEN_664;
  wire [31:0] _T_22 = ~_T_21;
  wire [10:0] lo_6 = {2'h0,reg_dcsr_cause,1'h0,2'h0,reg_dcsr_step,reg_dcsr_prv};
  wire [31:0] _T_23 = {4'h4,12'h0,reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku,1'h0,lo_6};
  wire [31:0] _T_24 = ~reg_dpc;
  wire [31:0] _T_27 = _T_24 | _GEN_664;
  wire [31:0] _T_28 = ~_T_27;
  wire [7:0] read_fcsr = {reg_frm,reg_fflags};
  wire [31:0] sie_mask = read_mideleg & 32'hefff;
  wire [31:0] read_sie = reg_mie & sie_mask;
  wire [31:0] read_sip = _GEN_41 & sie_mask;
  wire [8:0] lo_lo_6 = {io_status_spp,1'h0,1'h0,io_status_spie,1'h0,2'h0,io_status_sie,1'h0};
  wire [21:0] lo_7 = {2'h0,io_status_mxr,io_status_sum,1'h0,io_status_xs,io_status_fs,2'h0,io_status_vs,lo_lo_6};
  wire [104:0] _T_91 = {37'h0,4'h0,io_status_sd,23'h0,6'h0,io_status_uxl,io_status_sd_rv32,9'h0,lo_7};
  wire [31:0] _T_93 = {reg_satp_mode,9'h0,reg_satp_ppn};
  wire [31:0] _T_94 = ~reg_sepc;
  wire [31:0] _T_97 = _T_94 | _GEN_664;
  wire [31:0] _T_98 = ~_T_97;
  wire [7:0] _T_99 = {reg_pmp_0_cfg_l,2'h0,reg_pmp_0_cfg_a,reg_pmp_0_cfg_x,reg_pmp_0_cfg_w,reg_pmp_0_cfg_r};
  wire [7:0] _T_101 = {reg_pmp_2_cfg_l,2'h0,reg_pmp_2_cfg_a,reg_pmp_2_cfg_x,reg_pmp_2_cfg_w,reg_pmp_2_cfg_r};
  wire [15:0] lo_12 = {reg_pmp_1_cfg_l,2'h0,reg_pmp_1_cfg_a,reg_pmp_1_cfg_x,reg_pmp_1_cfg_w,reg_pmp_1_cfg_r,_T_99};
  wire [31:0] _T_103 = {reg_pmp_3_cfg_l,2'h0,reg_pmp_3_cfg_a,reg_pmp_3_cfg_x,reg_pmp_3_cfg_w,reg_pmp_3_cfg_r,_T_101,
    lo_12};
  wire [7:0] _T_104 = {reg_pmp_4_cfg_l,2'h0,reg_pmp_4_cfg_a,reg_pmp_4_cfg_x,reg_pmp_4_cfg_w,reg_pmp_4_cfg_r};
  wire [7:0] _T_106 = {reg_pmp_6_cfg_l,2'h0,reg_pmp_6_cfg_a,reg_pmp_6_cfg_x,reg_pmp_6_cfg_w,reg_pmp_6_cfg_r};
  wire [15:0] lo_17 = {reg_pmp_5_cfg_l,2'h0,reg_pmp_5_cfg_a,reg_pmp_5_cfg_x,reg_pmp_5_cfg_w,reg_pmp_5_cfg_r,_T_104};
  wire [31:0] _T_108 = {reg_pmp_7_cfg_l,2'h0,reg_pmp_7_cfg_a,reg_pmp_7_cfg_x,reg_pmp_7_cfg_w,reg_pmp_7_cfg_r,_T_106,
    lo_17};
  reg [31:0] reg_custom_0;
  wire [12:0] addr = {io_status_v,io_rw_addr};
  wire [11:0] decoded_decoded_plaInput = addr[11:0];
  wire [11:0] decoded_decoded_invInputs = ~decoded_decoded_plaInput;
  wire  decoded_decoded_andMatrixInput_0 = decoded_decoded_invInputs[1];
  wire  decoded_decoded_andMatrixInput_1 = decoded_decoded_invInputs[2];
  wire  decoded_decoded_andMatrixInput_2 = decoded_decoded_invInputs[3];
  wire  decoded_decoded_andMatrixInput_3 = decoded_decoded_invInputs[4];
  wire  decoded_decoded_andMatrixInput_4 = decoded_decoded_invInputs[5];
  wire  decoded_decoded_andMatrixInput_5 = decoded_decoded_invInputs[6];
  wire  decoded_decoded_andMatrixInput_6 = decoded_decoded_invInputs[7];
  wire  decoded_decoded_andMatrixInput_7 = decoded_decoded_invInputs[8];
  wire  decoded_decoded_andMatrixInput_8 = decoded_decoded_invInputs[9];
  wire  decoded_decoded_andMatrixInput_9 = decoded_decoded_invInputs[10];
  wire  decoded_decoded_andMatrixInput_10 = decoded_decoded_invInputs[11];
  wire [4:0] decoded_decoded_lo = {decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_7,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10};
  wire [10:0] _decoded_decoded_T = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo};
  wire  _decoded_decoded_T_1 = &_decoded_decoded_T;
  wire  decoded_decoded_andMatrixInput_0_1 = decoded_decoded_invInputs[0];
  wire  decoded_decoded_andMatrixInput_1_1 = decoded_decoded_plaInput[1];
  wire [5:0] decoded_decoded_lo_1 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10};
  wire [11:0] _decoded_decoded_T_2 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_1};
  wire  _decoded_decoded_T_3 = &_decoded_decoded_T_2;
  wire  decoded_decoded_andMatrixInput_0_2 = decoded_decoded_plaInput[0];
  wire [11:0] _decoded_decoded_T_4 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_1};
  wire  _decoded_decoded_T_5 = &_decoded_decoded_T_4;
  wire  decoded_decoded_andMatrixInput_6_3 = decoded_decoded_plaInput[8];
  wire [4:0] decoded_decoded_lo_3 = {decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10};
  wire [9:0] _decoded_decoded_T_6 = {decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10};
  wire  _decoded_decoded_T_7 = &_decoded_decoded_T_6;
  wire  decoded_decoded_andMatrixInput_2_4 = decoded_decoded_plaInput[2];
  wire [5:0] decoded_decoded_lo_4 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10};
  wire [11:0] _decoded_decoded_T_8 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_4};
  wire  _decoded_decoded_T_9 = &_decoded_decoded_T_8;
  wire [11:0] _decoded_decoded_T_10 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_4};
  wire  _decoded_decoded_T_11 = &_decoded_decoded_T_10;
  wire [10:0] _decoded_decoded_T_12 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_2_4,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_3};
  wire  _decoded_decoded_T_13 = &_decoded_decoded_T_12;
  wire  decoded_decoded_andMatrixInput_6_7 = decoded_decoded_plaInput[6];
  wire [5:0] decoded_decoded_lo_7 = {decoded_decoded_andMatrixInput_6_7,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10};
  wire [11:0] _decoded_decoded_T_14 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_7};
  wire  _decoded_decoded_T_15 = &_decoded_decoded_T_14;
  wire [11:0] _decoded_decoded_T_16 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_7};
  wire  _decoded_decoded_T_17 = &_decoded_decoded_T_16;
  wire [11:0] _decoded_decoded_T_18 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_7};
  wire  _decoded_decoded_T_19 = &_decoded_decoded_T_18;
  wire [11:0] _decoded_decoded_T_20 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_7};
  wire  _decoded_decoded_T_21 = &_decoded_decoded_T_20;
  wire [9:0] _decoded_decoded_T_22 = {decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_6_7,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10};
  wire  _decoded_decoded_T_23 = &_decoded_decoded_T_22;
  wire  decoded_decoded_andMatrixInput_0_12 = decoded_decoded_plaInput[7];
  wire [4:0] _decoded_decoded_T_24 = {decoded_decoded_andMatrixInput_0_12,decoded_decoded_andMatrixInput_6_3,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10};
  wire  _decoded_decoded_T_25 = &_decoded_decoded_T_24;
  wire  decoded_decoded_andMatrixInput_9_12 = decoded_decoded_plaInput[9];
  wire [5:0] decoded_decoded_lo_13 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10};
  wire [11:0] _decoded_decoded_T_26 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_27 = &_decoded_decoded_T_26;
  wire [11:0] _decoded_decoded_T_28 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_29 = &_decoded_decoded_T_28;
  wire [11:0] _decoded_decoded_T_30 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_31 = &_decoded_decoded_T_30;
  wire [11:0] _decoded_decoded_T_32 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_33 = &_decoded_decoded_T_32;
  wire [11:0] _decoded_decoded_T_34 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_35 = &_decoded_decoded_T_34;
  wire [11:0] _decoded_decoded_T_36 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_37 = &_decoded_decoded_T_36;
  wire [4:0] decoded_decoded_lo_19 = {decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,
    decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10};
  wire [10:0] _decoded_decoded_T_38 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_2_4,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_19};
  wire  _decoded_decoded_T_39 = &_decoded_decoded_T_38;
  wire  decoded_decoded_andMatrixInput_4_20 = decoded_decoded_plaInput[5];
  wire [10:0] _decoded_decoded_T_40 = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4_20,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_19};
  wire  _decoded_decoded_T_41 = &_decoded_decoded_T_40;
  wire [10:0] _decoded_decoded_T_42 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4_20,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_19};
  wire  _decoded_decoded_T_43 = &_decoded_decoded_T_42;
  wire [11:0] _decoded_decoded_T_44 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_45 = &_decoded_decoded_T_44;
  wire [11:0] _decoded_decoded_T_46 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_47 = &_decoded_decoded_T_46;
  wire [11:0] _decoded_decoded_T_48 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_49 = &_decoded_decoded_T_48;
  wire [11:0] _decoded_decoded_T_50 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_51 = &_decoded_decoded_T_50;
  wire  decoded_decoded_andMatrixInput_3_26 = decoded_decoded_plaInput[3];
  wire [11:0] _decoded_decoded_T_52 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_53 = &_decoded_decoded_T_52;
  wire [11:0] _decoded_decoded_T_54 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_55 = &_decoded_decoded_T_54;
  wire [11:0] _decoded_decoded_T_56 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_57 = &_decoded_decoded_T_56;
  wire [11:0] _decoded_decoded_T_58 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_59 = &_decoded_decoded_T_58;
  wire [11:0] _decoded_decoded_T_60 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_61 = &_decoded_decoded_T_60;
  wire [11:0] _decoded_decoded_T_62 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_63 = &_decoded_decoded_T_62;
  wire [11:0] _decoded_decoded_T_64 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_65 = &_decoded_decoded_T_64;
  wire [11:0] _decoded_decoded_T_66 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_67 = &_decoded_decoded_T_66;
  wire  decoded_decoded_andMatrixInput_4_34 = decoded_decoded_plaInput[4];
  wire [11:0] _decoded_decoded_T_68 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_69 = &_decoded_decoded_T_68;
  wire [11:0] _decoded_decoded_T_70 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_71 = &_decoded_decoded_T_70;
  wire [11:0] _decoded_decoded_T_72 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_73 = &_decoded_decoded_T_72;
  wire [11:0] _decoded_decoded_T_74 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_75 = &_decoded_decoded_T_74;
  wire [11:0] _decoded_decoded_T_76 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_77 = &_decoded_decoded_T_76;
  wire [11:0] _decoded_decoded_T_78 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_79 = &_decoded_decoded_T_78;
  wire [11:0] _decoded_decoded_T_80 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_81 = &_decoded_decoded_T_80;
  wire [11:0] _decoded_decoded_T_82 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_83 = &_decoded_decoded_T_82;
  wire [11:0] _decoded_decoded_T_84 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_85 = &_decoded_decoded_T_84;
  wire [11:0] _decoded_decoded_T_86 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_87 = &_decoded_decoded_T_86;
  wire [11:0] _decoded_decoded_T_88 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_89 = &_decoded_decoded_T_88;
  wire [11:0] _decoded_decoded_T_90 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_91 = &_decoded_decoded_T_90;
  wire [11:0] _decoded_decoded_T_92 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_93 = &_decoded_decoded_T_92;
  wire [11:0] _decoded_decoded_T_94 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_95 = &_decoded_decoded_T_94;
  wire [11:0] _decoded_decoded_T_96 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_97 = &_decoded_decoded_T_96;
  wire [11:0] _decoded_decoded_T_98 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_13};
  wire  _decoded_decoded_T_99 = &_decoded_decoded_T_98;
  wire [5:0] decoded_decoded_lo_50 = {decoded_decoded_andMatrixInput_6_7,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10};
  wire [11:0] _decoded_decoded_T_100 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_50};
  wire  _decoded_decoded_T_101 = &_decoded_decoded_T_100;
  wire [11:0] _decoded_decoded_T_102 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_50};
  wire  _decoded_decoded_T_103 = &_decoded_decoded_T_102;
  wire [11:0] _decoded_decoded_T_104 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_50};
  wire  _decoded_decoded_T_105 = &_decoded_decoded_T_104;
  wire [11:0] _decoded_decoded_T_106 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_50};
  wire  _decoded_decoded_T_107 = &_decoded_decoded_T_106;
  wire [9:0] _decoded_decoded_T_108 = {decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_6_7,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,
    decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10};
  wire  _decoded_decoded_T_109 = &_decoded_decoded_T_108;
  wire [5:0] decoded_decoded_lo_55 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_0_12,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10};
  wire [11:0] _decoded_decoded_T_110 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_111 = &_decoded_decoded_T_110;
  wire [11:0] _decoded_decoded_T_112 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_113 = &_decoded_decoded_T_112;
  wire [11:0] _decoded_decoded_T_114 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_115 = &_decoded_decoded_T_114;
  wire [11:0] _decoded_decoded_T_116 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_117 = &_decoded_decoded_T_116;
  wire [11:0] _decoded_decoded_T_118 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_119 = &_decoded_decoded_T_118;
  wire [11:0] _decoded_decoded_T_120 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_121 = &_decoded_decoded_T_120;
  wire [11:0] _decoded_decoded_T_122 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_123 = &_decoded_decoded_T_122;
  wire [11:0] _decoded_decoded_T_124 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_125 = &_decoded_decoded_T_124;
  wire [11:0] _decoded_decoded_T_126 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_127 = &_decoded_decoded_T_126;
  wire [11:0] _decoded_decoded_T_128 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_129 = &_decoded_decoded_T_128;
  wire [11:0] _decoded_decoded_T_130 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_131 = &_decoded_decoded_T_130;
  wire [11:0] _decoded_decoded_T_132 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_133 = &_decoded_decoded_T_132;
  wire [11:0] _decoded_decoded_T_134 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_135 = &_decoded_decoded_T_134;
  wire [11:0] _decoded_decoded_T_136 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_137 = &_decoded_decoded_T_136;
  wire [11:0] _decoded_decoded_T_138 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_139 = &_decoded_decoded_T_138;
  wire [11:0] _decoded_decoded_T_140 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_141 = &_decoded_decoded_T_140;
  wire [11:0] _decoded_decoded_T_142 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_143 = &_decoded_decoded_T_142;
  wire [11:0] _decoded_decoded_T_144 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_145 = &_decoded_decoded_T_144;
  wire [11:0] _decoded_decoded_T_146 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_147 = &_decoded_decoded_T_146;
  wire [11:0] _decoded_decoded_T_148 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_55};
  wire  _decoded_decoded_T_149 = &_decoded_decoded_T_148;
  wire  decoded_decoded_andMatrixInput_10_71 = decoded_decoded_plaInput[10];
  wire [5:0] decoded_decoded_lo_75 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_0_12,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_10_71,
    decoded_decoded_andMatrixInput_10};
  wire [11:0] _decoded_decoded_T_150 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_75};
  wire  _decoded_decoded_T_151 = &_decoded_decoded_T_150;
  wire [11:0] _decoded_decoded_T_152 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_75};
  wire  _decoded_decoded_T_153 = &_decoded_decoded_T_152;
  wire [11:0] _decoded_decoded_T_154 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_75};
  wire  _decoded_decoded_T_155 = &_decoded_decoded_T_154;
  wire [11:0] _decoded_decoded_T_156 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_75};
  wire  _decoded_decoded_T_157 = &_decoded_decoded_T_156;
  wire [11:0] _decoded_decoded_T_158 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_75};
  wire  _decoded_decoded_T_159 = &_decoded_decoded_T_158;
  wire [11:0] _decoded_decoded_T_160 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4_20,decoded_decoded_lo_75};
  wire  _decoded_decoded_T_161 = &_decoded_decoded_T_160;
  wire [4:0] decoded_decoded_lo_81 = {decoded_decoded_andMatrixInput_0_12,decoded_decoded_andMatrixInput_6_3,
    decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_10_71,decoded_decoded_andMatrixInput_10};
  wire [10:0] _decoded_decoded_T_162 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,decoded_decoded_andMatrixInput_4_20,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_81};
  wire  _decoded_decoded_T_163 = &_decoded_decoded_T_162;
  wire [5:0] _decoded_decoded_T_164 = {decoded_decoded_andMatrixInput_6_7,decoded_decoded_andMatrixInput_0_12,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_10_71,
    decoded_decoded_andMatrixInput_10};
  wire  _decoded_decoded_T_165 = &_decoded_decoded_T_164;
  wire  decoded_decoded_andMatrixInput_10_78 = decoded_decoded_plaInput[11];
  wire [4:0] decoded_decoded_lo_83 = {decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,
    decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10_78};
  wire [10:0] _decoded_decoded_T_166 = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_83};
  wire  _decoded_decoded_T_167 = &_decoded_decoded_T_166;
  wire [5:0] decoded_decoded_lo_84 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10_78};
  wire [11:0] _decoded_decoded_T_168 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_169 = &_decoded_decoded_T_168;
  wire [11:0] _decoded_decoded_T_170 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_171 = &_decoded_decoded_T_170;
  wire [11:0] _decoded_decoded_T_172 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_173 = &_decoded_decoded_T_172;
  wire [11:0] _decoded_decoded_T_174 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_175 = &_decoded_decoded_T_174;
  wire [11:0] _decoded_decoded_T_176 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_177 = &_decoded_decoded_T_176;
  wire [11:0] _decoded_decoded_T_178 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_179 = &_decoded_decoded_T_178;
  wire [11:0] _decoded_decoded_T_180 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_181 = &_decoded_decoded_T_180;
  wire [11:0] _decoded_decoded_T_182 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_183 = &_decoded_decoded_T_182;
  wire [11:0] _decoded_decoded_T_184 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_185 = &_decoded_decoded_T_184;
  wire [11:0] _decoded_decoded_T_186 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_187 = &_decoded_decoded_T_186;
  wire [11:0] _decoded_decoded_T_188 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_189 = &_decoded_decoded_T_188;
  wire [11:0] _decoded_decoded_T_190 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_191 = &_decoded_decoded_T_190;
  wire [11:0] _decoded_decoded_T_192 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_193 = &_decoded_decoded_T_192;
  wire [11:0] _decoded_decoded_T_194 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_195 = &_decoded_decoded_T_194;
  wire [11:0] _decoded_decoded_T_196 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_197 = &_decoded_decoded_T_196;
  wire [11:0] _decoded_decoded_T_198 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_199 = &_decoded_decoded_T_198;
  wire [11:0] _decoded_decoded_T_200 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_201 = &_decoded_decoded_T_200;
  wire [11:0] _decoded_decoded_T_202 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_203 = &_decoded_decoded_T_202;
  wire [11:0] _decoded_decoded_T_204 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_205 = &_decoded_decoded_T_204;
  wire [11:0] _decoded_decoded_T_206 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_207 = &_decoded_decoded_T_206;
  wire [11:0] _decoded_decoded_T_208 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_209 = &_decoded_decoded_T_208;
  wire [11:0] _decoded_decoded_T_210 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_211 = &_decoded_decoded_T_210;
  wire [11:0] _decoded_decoded_T_212 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_213 = &_decoded_decoded_T_212;
  wire [11:0] _decoded_decoded_T_214 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_215 = &_decoded_decoded_T_214;
  wire [11:0] _decoded_decoded_T_216 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_217 = &_decoded_decoded_T_216;
  wire [11:0] _decoded_decoded_T_218 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_219 = &_decoded_decoded_T_218;
  wire [11:0] _decoded_decoded_T_220 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_221 = &_decoded_decoded_T_220;
  wire [11:0] _decoded_decoded_T_222 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_223 = &_decoded_decoded_T_222;
  wire [11:0] _decoded_decoded_T_224 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_225 = &_decoded_decoded_T_224;
  wire [11:0] _decoded_decoded_T_226 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_84};
  wire  _decoded_decoded_T_227 = &_decoded_decoded_T_226;
  wire [4:0] decoded_decoded_lo_114 = {decoded_decoded_andMatrixInput_0_12,decoded_decoded_andMatrixInput_6_3,
    decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,decoded_decoded_andMatrixInput_10_78};
  wire [10:0] _decoded_decoded_T_228 = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_114};
  wire  _decoded_decoded_T_229 = &_decoded_decoded_T_228;
  wire [5:0] decoded_decoded_lo_115 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_0_12,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_9,
    decoded_decoded_andMatrixInput_10_78};
  wire [11:0] _decoded_decoded_T_230 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_231 = &_decoded_decoded_T_230;
  wire [11:0] _decoded_decoded_T_232 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_233 = &_decoded_decoded_T_232;
  wire [11:0] _decoded_decoded_T_234 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_235 = &_decoded_decoded_T_234;
  wire [11:0] _decoded_decoded_T_236 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_237 = &_decoded_decoded_T_236;
  wire [11:0] _decoded_decoded_T_238 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_239 = &_decoded_decoded_T_238;
  wire [11:0] _decoded_decoded_T_240 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_241 = &_decoded_decoded_T_240;
  wire [11:0] _decoded_decoded_T_242 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_243 = &_decoded_decoded_T_242;
  wire [11:0] _decoded_decoded_T_244 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_245 = &_decoded_decoded_T_244;
  wire [11:0] _decoded_decoded_T_246 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_247 = &_decoded_decoded_T_246;
  wire [11:0] _decoded_decoded_T_248 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_249 = &_decoded_decoded_T_248;
  wire [11:0] _decoded_decoded_T_250 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_251 = &_decoded_decoded_T_250;
  wire [11:0] _decoded_decoded_T_252 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_253 = &_decoded_decoded_T_252;
  wire [11:0] _decoded_decoded_T_254 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_255 = &_decoded_decoded_T_254;
  wire [11:0] _decoded_decoded_T_256 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_257 = &_decoded_decoded_T_256;
  wire [11:0] _decoded_decoded_T_258 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_259 = &_decoded_decoded_T_258;
  wire [11:0] _decoded_decoded_T_260 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_261 = &_decoded_decoded_T_260;
  wire [11:0] _decoded_decoded_T_262 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_263 = &_decoded_decoded_T_262;
  wire [11:0] _decoded_decoded_T_264 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_265 = &_decoded_decoded_T_264;
  wire [11:0] _decoded_decoded_T_266 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_267 = &_decoded_decoded_T_266;
  wire [11:0] _decoded_decoded_T_268 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_269 = &_decoded_decoded_T_268;
  wire [11:0] _decoded_decoded_T_270 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_271 = &_decoded_decoded_T_270;
  wire [11:0] _decoded_decoded_T_272 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_273 = &_decoded_decoded_T_272;
  wire [11:0] _decoded_decoded_T_274 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_275 = &_decoded_decoded_T_274;
  wire [11:0] _decoded_decoded_T_276 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_277 = &_decoded_decoded_T_276;
  wire [11:0] _decoded_decoded_T_278 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_279 = &_decoded_decoded_T_278;
  wire [11:0] _decoded_decoded_T_280 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_281 = &_decoded_decoded_T_280;
  wire [11:0] _decoded_decoded_T_282 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_283 = &_decoded_decoded_T_282;
  wire [11:0] _decoded_decoded_T_284 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_285 = &_decoded_decoded_T_284;
  wire [11:0] _decoded_decoded_T_286 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_287 = &_decoded_decoded_T_286;
  wire [11:0] _decoded_decoded_T_288 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_115};
  wire  _decoded_decoded_T_289 = &_decoded_decoded_T_288;
  wire [4:0] decoded_decoded_lo_145 = {decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_7,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_10_71,decoded_decoded_andMatrixInput_10_78};
  wire [10:0] _decoded_decoded_T_290 = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_145};
  wire  _decoded_decoded_T_291 = &_decoded_decoded_T_290;
  wire [5:0] decoded_decoded_lo_146 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_10_71,
    decoded_decoded_andMatrixInput_10_78};
  wire [11:0] _decoded_decoded_T_292 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_293 = &_decoded_decoded_T_292;
  wire [11:0] _decoded_decoded_T_294 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_295 = &_decoded_decoded_T_294;
  wire [11:0] _decoded_decoded_T_296 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_297 = &_decoded_decoded_T_296;
  wire [11:0] _decoded_decoded_T_298 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_299 = &_decoded_decoded_T_298;
  wire [11:0] _decoded_decoded_T_300 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_301 = &_decoded_decoded_T_300;
  wire [11:0] _decoded_decoded_T_302 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_303 = &_decoded_decoded_T_302;
  wire [11:0] _decoded_decoded_T_304 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_305 = &_decoded_decoded_T_304;
  wire [11:0] _decoded_decoded_T_306 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_307 = &_decoded_decoded_T_306;
  wire [11:0] _decoded_decoded_T_308 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_309 = &_decoded_decoded_T_308;
  wire [11:0] _decoded_decoded_T_310 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_311 = &_decoded_decoded_T_310;
  wire [11:0] _decoded_decoded_T_312 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_313 = &_decoded_decoded_T_312;
  wire [11:0] _decoded_decoded_T_314 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_315 = &_decoded_decoded_T_314;
  wire [11:0] _decoded_decoded_T_316 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_317 = &_decoded_decoded_T_316;
  wire [11:0] _decoded_decoded_T_318 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_319 = &_decoded_decoded_T_318;
  wire [11:0] _decoded_decoded_T_320 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_321 = &_decoded_decoded_T_320;
  wire [11:0] _decoded_decoded_T_322 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_323 = &_decoded_decoded_T_322;
  wire [11:0] _decoded_decoded_T_324 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_325 = &_decoded_decoded_T_324;
  wire [11:0] _decoded_decoded_T_326 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_327 = &_decoded_decoded_T_326;
  wire [11:0] _decoded_decoded_T_328 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_329 = &_decoded_decoded_T_328;
  wire [11:0] _decoded_decoded_T_330 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_331 = &_decoded_decoded_T_330;
  wire [11:0] _decoded_decoded_T_332 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_333 = &_decoded_decoded_T_332;
  wire [11:0] _decoded_decoded_T_334 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_335 = &_decoded_decoded_T_334;
  wire [11:0] _decoded_decoded_T_336 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_337 = &_decoded_decoded_T_336;
  wire [11:0] _decoded_decoded_T_338 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_339 = &_decoded_decoded_T_338;
  wire [11:0] _decoded_decoded_T_340 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_341 = &_decoded_decoded_T_340;
  wire [11:0] _decoded_decoded_T_342 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_343 = &_decoded_decoded_T_342;
  wire [11:0] _decoded_decoded_T_344 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_345 = &_decoded_decoded_T_344;
  wire [11:0] _decoded_decoded_T_346 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_347 = &_decoded_decoded_T_346;
  wire [11:0] _decoded_decoded_T_348 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_349 = &_decoded_decoded_T_348;
  wire [11:0] _decoded_decoded_T_350 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_146};
  wire  _decoded_decoded_T_351 = &_decoded_decoded_T_350;
  wire [4:0] decoded_decoded_lo_176 = {decoded_decoded_andMatrixInput_0_12,decoded_decoded_andMatrixInput_7,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_10_71,decoded_decoded_andMatrixInput_10_78};
  wire [10:0] _decoded_decoded_T_352 = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_176};
  wire  _decoded_decoded_T_353 = &_decoded_decoded_T_352;
  wire [5:0] decoded_decoded_lo_177 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_0_12,
    decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_10_71,
    decoded_decoded_andMatrixInput_10_78};
  wire [11:0] _decoded_decoded_T_354 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_355 = &_decoded_decoded_T_354;
  wire [11:0] _decoded_decoded_T_356 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_357 = &_decoded_decoded_T_356;
  wire [11:0] _decoded_decoded_T_358 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_359 = &_decoded_decoded_T_358;
  wire [11:0] _decoded_decoded_T_360 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_361 = &_decoded_decoded_T_360;
  wire [11:0] _decoded_decoded_T_362 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_363 = &_decoded_decoded_T_362;
  wire [11:0] _decoded_decoded_T_364 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_365 = &_decoded_decoded_T_364;
  wire [11:0] _decoded_decoded_T_366 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_367 = &_decoded_decoded_T_366;
  wire [11:0] _decoded_decoded_T_368 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_369 = &_decoded_decoded_T_368;
  wire [11:0] _decoded_decoded_T_370 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_371 = &_decoded_decoded_T_370;
  wire [11:0] _decoded_decoded_T_372 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_373 = &_decoded_decoded_T_372;
  wire [11:0] _decoded_decoded_T_374 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_375 = &_decoded_decoded_T_374;
  wire [11:0] _decoded_decoded_T_376 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_377 = &_decoded_decoded_T_376;
  wire [11:0] _decoded_decoded_T_378 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_379 = &_decoded_decoded_T_378;
  wire [11:0] _decoded_decoded_T_380 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_381 = &_decoded_decoded_T_380;
  wire [11:0] _decoded_decoded_T_382 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_383 = &_decoded_decoded_T_382;
  wire [11:0] _decoded_decoded_T_384 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_385 = &_decoded_decoded_T_384;
  wire [11:0] _decoded_decoded_T_386 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_387 = &_decoded_decoded_T_386;
  wire [11:0] _decoded_decoded_T_388 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_389 = &_decoded_decoded_T_388;
  wire [11:0] _decoded_decoded_T_390 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_391 = &_decoded_decoded_T_390;
  wire [11:0] _decoded_decoded_T_392 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_393 = &_decoded_decoded_T_392;
  wire [11:0] _decoded_decoded_T_394 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_395 = &_decoded_decoded_T_394;
  wire [11:0] _decoded_decoded_T_396 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_397 = &_decoded_decoded_T_396;
  wire [11:0] _decoded_decoded_T_398 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_399 = &_decoded_decoded_T_398;
  wire [11:0] _decoded_decoded_T_400 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_401 = &_decoded_decoded_T_400;
  wire [11:0] _decoded_decoded_T_402 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_403 = &_decoded_decoded_T_402;
  wire [11:0] _decoded_decoded_T_404 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_405 = &_decoded_decoded_T_404;
  wire [11:0] _decoded_decoded_T_406 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_407 = &_decoded_decoded_T_406;
  wire [11:0] _decoded_decoded_T_408 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_409 = &_decoded_decoded_T_408;
  wire [11:0] _decoded_decoded_T_410 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_411 = &_decoded_decoded_T_410;
  wire [11:0] _decoded_decoded_T_412 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_3_26,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_177};
  wire  _decoded_decoded_T_413 = &_decoded_decoded_T_412;
  wire [4:0] decoded_decoded_lo_207 = {decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,
    decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_10_71,decoded_decoded_andMatrixInput_10_78};
  wire [10:0] _decoded_decoded_T_414 = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_lo_207};
  wire  _decoded_decoded_T_415 = &_decoded_decoded_T_414;
  wire [5:0] decoded_decoded_lo_208 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,decoded_decoded_andMatrixInput_10_71,
    decoded_decoded_andMatrixInput_10_78};
  wire [11:0] _decoded_decoded_T_416 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_208};
  wire  _decoded_decoded_T_417 = &_decoded_decoded_T_416;
  wire [11:0] _decoded_decoded_T_418 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_34,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_208};
  wire  _decoded_decoded_T_419 = &_decoded_decoded_T_418;
  wire [9:0] _decoded_decoded_T_420 = {decoded_decoded_andMatrixInput_2_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_34,decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_6_3,decoded_decoded_andMatrixInput_9_12,
    decoded_decoded_andMatrixInput_10_71,decoded_decoded_andMatrixInput_10_78};
  wire  _decoded_decoded_T_421 = &_decoded_decoded_T_420;
  wire  _decoded_decoded_orMatrixOutputs_T = |_decoded_decoded_T_419;
  wire  _decoded_decoded_orMatrixOutputs_T_1 = |_decoded_decoded_T_415;
  wire  _decoded_decoded_orMatrixOutputs_T_2 = |_decoded_decoded_T_417;
  wire  _decoded_decoded_orMatrixOutputs_T_3 = |_decoded_decoded_T_165;
  wire  _decoded_decoded_orMatrixOutputs_T_4 = |_decoded_decoded_T_149;
  wire  _decoded_decoded_orMatrixOutputs_T_5 = |_decoded_decoded_T_147;
  wire  _decoded_decoded_orMatrixOutputs_T_6 = |_decoded_decoded_T_145;
  wire  _decoded_decoded_orMatrixOutputs_T_7 = |_decoded_decoded_T_143;
  wire  _decoded_decoded_orMatrixOutputs_T_8 = |_decoded_decoded_T_141;
  wire  _decoded_decoded_orMatrixOutputs_T_9 = |_decoded_decoded_T_139;
  wire  _decoded_decoded_orMatrixOutputs_T_10 = |_decoded_decoded_T_137;
  wire  _decoded_decoded_orMatrixOutputs_T_11 = |_decoded_decoded_T_135;
  wire  _decoded_decoded_orMatrixOutputs_T_12 = |_decoded_decoded_T_133;
  wire  _decoded_decoded_orMatrixOutputs_T_13 = |_decoded_decoded_T_131;
  wire  _decoded_decoded_orMatrixOutputs_T_14 = |_decoded_decoded_T_129;
  wire  _decoded_decoded_orMatrixOutputs_T_15 = |_decoded_decoded_T_127;
  wire  _decoded_decoded_orMatrixOutputs_T_16 = |_decoded_decoded_T_125;
  wire  _decoded_decoded_orMatrixOutputs_T_17 = |_decoded_decoded_T_123;
  wire  _decoded_decoded_orMatrixOutputs_T_18 = |_decoded_decoded_T_121;
  wire  _decoded_decoded_orMatrixOutputs_T_19 = |_decoded_decoded_T_119;
  wire  _decoded_decoded_orMatrixOutputs_T_20 = |_decoded_decoded_T_117;
  wire  _decoded_decoded_orMatrixOutputs_T_21 = |_decoded_decoded_T_115;
  wire  _decoded_decoded_orMatrixOutputs_T_22 = |_decoded_decoded_T_113;
  wire  _decoded_decoded_orMatrixOutputs_T_23 = |_decoded_decoded_T_111;
  wire  _decoded_decoded_orMatrixOutputs_T_24 = |_decoded_decoded_T_31;
  wire  _decoded_decoded_orMatrixOutputs_T_25 = |_decoded_decoded_T_33;
  wire  _decoded_decoded_orMatrixOutputs_T_26 = |_decoded_decoded_T_13;
  wire  _decoded_decoded_orMatrixOutputs_T_27 = |_decoded_decoded_T_11;
  wire  _decoded_decoded_orMatrixOutputs_T_28 = |_decoded_decoded_T_17;
  wire  _decoded_decoded_orMatrixOutputs_T_29 = |_decoded_decoded_T_25;
  wire  _decoded_decoded_orMatrixOutputs_T_30 = |_decoded_decoded_T_21;
  wire  _decoded_decoded_orMatrixOutputs_T_31 = |_decoded_decoded_T_19;
  wire  _decoded_decoded_orMatrixOutputs_T_32 = |_decoded_decoded_T_15;
  wire  _decoded_decoded_orMatrixOutputs_T_33 = |_decoded_decoded_T_9;
  wire  _decoded_decoded_orMatrixOutputs_T_34 = |_decoded_decoded_T_23;
  wire  _decoded_decoded_orMatrixOutputs_T_35 = |_decoded_decoded_T_7;
  wire  _decoded_decoded_orMatrixOutputs_T_36 = |_decoded_decoded_T_355;
  wire  _decoded_decoded_orMatrixOutputs_T_37 = |_decoded_decoded_T_353;
  wire  _decoded_decoded_orMatrixOutputs_T_38 = |_decoded_decoded_T_231;
  wire  _decoded_decoded_orMatrixOutputs_T_39 = |_decoded_decoded_T_229;
  wire  _decoded_decoded_orMatrixOutputs_T_40 = |_decoded_decoded_T_293;
  wire  _decoded_decoded_orMatrixOutputs_T_41 = |_decoded_decoded_T_291;
  wire  _decoded_decoded_orMatrixOutputs_T_42 = |_decoded_decoded_T_39;
  wire  _decoded_decoded_orMatrixOutputs_T_43 = |_decoded_decoded_T_413;
  wire  _decoded_decoded_orMatrixOutputs_T_44 = |_decoded_decoded_T_289;
  wire  _decoded_decoded_orMatrixOutputs_T_45 = |_decoded_decoded_T_351;
  wire  _decoded_decoded_orMatrixOutputs_T_46 = |_decoded_decoded_T_227;
  wire  _decoded_decoded_orMatrixOutputs_T_47 = |_decoded_decoded_T_99;
  wire  _decoded_decoded_orMatrixOutputs_T_48 = |_decoded_decoded_T_411;
  wire  _decoded_decoded_orMatrixOutputs_T_49 = |_decoded_decoded_T_287;
  wire  _decoded_decoded_orMatrixOutputs_T_50 = |_decoded_decoded_T_349;
  wire  _decoded_decoded_orMatrixOutputs_T_51 = |_decoded_decoded_T_225;
  wire  _decoded_decoded_orMatrixOutputs_T_52 = |_decoded_decoded_T_97;
  wire  _decoded_decoded_orMatrixOutputs_T_53 = |_decoded_decoded_T_409;
  wire  _decoded_decoded_orMatrixOutputs_T_54 = |_decoded_decoded_T_285;
  wire  _decoded_decoded_orMatrixOutputs_T_55 = |_decoded_decoded_T_347;
  wire  _decoded_decoded_orMatrixOutputs_T_56 = |_decoded_decoded_T_223;
  wire  _decoded_decoded_orMatrixOutputs_T_57 = |_decoded_decoded_T_95;
  wire  _decoded_decoded_orMatrixOutputs_T_58 = |_decoded_decoded_T_407;
  wire  _decoded_decoded_orMatrixOutputs_T_59 = |_decoded_decoded_T_283;
  wire  _decoded_decoded_orMatrixOutputs_T_60 = |_decoded_decoded_T_345;
  wire  _decoded_decoded_orMatrixOutputs_T_61 = |_decoded_decoded_T_221;
  wire  _decoded_decoded_orMatrixOutputs_T_62 = |_decoded_decoded_T_93;
  wire  _decoded_decoded_orMatrixOutputs_T_63 = |_decoded_decoded_T_405;
  wire  _decoded_decoded_orMatrixOutputs_T_64 = |_decoded_decoded_T_281;
  wire  _decoded_decoded_orMatrixOutputs_T_65 = |_decoded_decoded_T_343;
  wire  _decoded_decoded_orMatrixOutputs_T_66 = |_decoded_decoded_T_219;
  wire  _decoded_decoded_orMatrixOutputs_T_67 = |_decoded_decoded_T_91;
  wire  _decoded_decoded_orMatrixOutputs_T_68 = |_decoded_decoded_T_403;
  wire  _decoded_decoded_orMatrixOutputs_T_69 = |_decoded_decoded_T_279;
  wire  _decoded_decoded_orMatrixOutputs_T_70 = |_decoded_decoded_T_341;
  wire  _decoded_decoded_orMatrixOutputs_T_71 = |_decoded_decoded_T_217;
  wire  _decoded_decoded_orMatrixOutputs_T_72 = |_decoded_decoded_T_89;
  wire  _decoded_decoded_orMatrixOutputs_T_73 = |_decoded_decoded_T_401;
  wire  _decoded_decoded_orMatrixOutputs_T_74 = |_decoded_decoded_T_277;
  wire  _decoded_decoded_orMatrixOutputs_T_75 = |_decoded_decoded_T_339;
  wire  _decoded_decoded_orMatrixOutputs_T_76 = |_decoded_decoded_T_215;
  wire  _decoded_decoded_orMatrixOutputs_T_77 = |_decoded_decoded_T_87;
  wire  _decoded_decoded_orMatrixOutputs_T_78 = |_decoded_decoded_T_399;
  wire  _decoded_decoded_orMatrixOutputs_T_79 = |_decoded_decoded_T_275;
  wire  _decoded_decoded_orMatrixOutputs_T_80 = |_decoded_decoded_T_337;
  wire  _decoded_decoded_orMatrixOutputs_T_81 = |_decoded_decoded_T_213;
  wire  _decoded_decoded_orMatrixOutputs_T_82 = |_decoded_decoded_T_85;
  wire  _decoded_decoded_orMatrixOutputs_T_83 = |_decoded_decoded_T_397;
  wire  _decoded_decoded_orMatrixOutputs_T_84 = |_decoded_decoded_T_273;
  wire  _decoded_decoded_orMatrixOutputs_T_85 = |_decoded_decoded_T_335;
  wire  _decoded_decoded_orMatrixOutputs_T_86 = |_decoded_decoded_T_211;
  wire  _decoded_decoded_orMatrixOutputs_T_87 = |_decoded_decoded_T_83;
  wire  _decoded_decoded_orMatrixOutputs_T_88 = |_decoded_decoded_T_395;
  wire  _decoded_decoded_orMatrixOutputs_T_89 = |_decoded_decoded_T_271;
  wire  _decoded_decoded_orMatrixOutputs_T_90 = |_decoded_decoded_T_333;
  wire  _decoded_decoded_orMatrixOutputs_T_91 = |_decoded_decoded_T_209;
  wire  _decoded_decoded_orMatrixOutputs_T_92 = |_decoded_decoded_T_81;
  wire  _decoded_decoded_orMatrixOutputs_T_93 = |_decoded_decoded_T_393;
  wire  _decoded_decoded_orMatrixOutputs_T_94 = |_decoded_decoded_T_269;
  wire  _decoded_decoded_orMatrixOutputs_T_95 = |_decoded_decoded_T_331;
  wire  _decoded_decoded_orMatrixOutputs_T_96 = |_decoded_decoded_T_207;
  wire  _decoded_decoded_orMatrixOutputs_T_97 = |_decoded_decoded_T_79;
  wire  _decoded_decoded_orMatrixOutputs_T_98 = |_decoded_decoded_T_391;
  wire  _decoded_decoded_orMatrixOutputs_T_99 = |_decoded_decoded_T_267;
  wire  _decoded_decoded_orMatrixOutputs_T_100 = |_decoded_decoded_T_329;
  wire  _decoded_decoded_orMatrixOutputs_T_101 = |_decoded_decoded_T_205;
  wire  _decoded_decoded_orMatrixOutputs_T_102 = |_decoded_decoded_T_77;
  wire  _decoded_decoded_orMatrixOutputs_T_103 = |_decoded_decoded_T_389;
  wire  _decoded_decoded_orMatrixOutputs_T_104 = |_decoded_decoded_T_265;
  wire  _decoded_decoded_orMatrixOutputs_T_105 = |_decoded_decoded_T_327;
  wire  _decoded_decoded_orMatrixOutputs_T_106 = |_decoded_decoded_T_203;
  wire  _decoded_decoded_orMatrixOutputs_T_107 = |_decoded_decoded_T_75;
  wire  _decoded_decoded_orMatrixOutputs_T_108 = |_decoded_decoded_T_387;
  wire  _decoded_decoded_orMatrixOutputs_T_109 = |_decoded_decoded_T_263;
  wire  _decoded_decoded_orMatrixOutputs_T_110 = |_decoded_decoded_T_325;
  wire  _decoded_decoded_orMatrixOutputs_T_111 = |_decoded_decoded_T_201;
  wire  _decoded_decoded_orMatrixOutputs_T_112 = |_decoded_decoded_T_73;
  wire  _decoded_decoded_orMatrixOutputs_T_113 = |_decoded_decoded_T_385;
  wire  _decoded_decoded_orMatrixOutputs_T_114 = |_decoded_decoded_T_261;
  wire  _decoded_decoded_orMatrixOutputs_T_115 = |_decoded_decoded_T_323;
  wire  _decoded_decoded_orMatrixOutputs_T_116 = |_decoded_decoded_T_199;
  wire  _decoded_decoded_orMatrixOutputs_T_117 = |_decoded_decoded_T_71;
  wire  _decoded_decoded_orMatrixOutputs_T_118 = |_decoded_decoded_T_383;
  wire  _decoded_decoded_orMatrixOutputs_T_119 = |_decoded_decoded_T_259;
  wire  _decoded_decoded_orMatrixOutputs_T_120 = |_decoded_decoded_T_321;
  wire  _decoded_decoded_orMatrixOutputs_T_121 = |_decoded_decoded_T_197;
  wire  _decoded_decoded_orMatrixOutputs_T_122 = |_decoded_decoded_T_69;
  wire  _decoded_decoded_orMatrixOutputs_T_123 = |_decoded_decoded_T_381;
  wire  _decoded_decoded_orMatrixOutputs_T_124 = |_decoded_decoded_T_257;
  wire  _decoded_decoded_orMatrixOutputs_T_125 = |_decoded_decoded_T_319;
  wire  _decoded_decoded_orMatrixOutputs_T_126 = |_decoded_decoded_T_195;
  wire  _decoded_decoded_orMatrixOutputs_T_127 = |_decoded_decoded_T_67;
  wire  _decoded_decoded_orMatrixOutputs_T_128 = |_decoded_decoded_T_379;
  wire  _decoded_decoded_orMatrixOutputs_T_129 = |_decoded_decoded_T_255;
  wire  _decoded_decoded_orMatrixOutputs_T_130 = |_decoded_decoded_T_317;
  wire  _decoded_decoded_orMatrixOutputs_T_131 = |_decoded_decoded_T_193;
  wire  _decoded_decoded_orMatrixOutputs_T_132 = |_decoded_decoded_T_65;
  wire  _decoded_decoded_orMatrixOutputs_T_133 = |_decoded_decoded_T_377;
  wire  _decoded_decoded_orMatrixOutputs_T_134 = |_decoded_decoded_T_253;
  wire  _decoded_decoded_orMatrixOutputs_T_135 = |_decoded_decoded_T_315;
  wire  _decoded_decoded_orMatrixOutputs_T_136 = |_decoded_decoded_T_191;
  wire  _decoded_decoded_orMatrixOutputs_T_137 = |_decoded_decoded_T_63;
  wire  _decoded_decoded_orMatrixOutputs_T_138 = |_decoded_decoded_T_375;
  wire  _decoded_decoded_orMatrixOutputs_T_139 = |_decoded_decoded_T_251;
  wire  _decoded_decoded_orMatrixOutputs_T_140 = |_decoded_decoded_T_313;
  wire  _decoded_decoded_orMatrixOutputs_T_141 = |_decoded_decoded_T_189;
  wire  _decoded_decoded_orMatrixOutputs_T_142 = |_decoded_decoded_T_61;
  wire  _decoded_decoded_orMatrixOutputs_T_143 = |_decoded_decoded_T_373;
  wire  _decoded_decoded_orMatrixOutputs_T_144 = |_decoded_decoded_T_249;
  wire  _decoded_decoded_orMatrixOutputs_T_145 = |_decoded_decoded_T_311;
  wire  _decoded_decoded_orMatrixOutputs_T_146 = |_decoded_decoded_T_187;
  wire  _decoded_decoded_orMatrixOutputs_T_147 = |_decoded_decoded_T_59;
  wire  _decoded_decoded_orMatrixOutputs_T_148 = |_decoded_decoded_T_371;
  wire  _decoded_decoded_orMatrixOutputs_T_149 = |_decoded_decoded_T_247;
  wire  _decoded_decoded_orMatrixOutputs_T_150 = |_decoded_decoded_T_309;
  wire  _decoded_decoded_orMatrixOutputs_T_151 = |_decoded_decoded_T_185;
  wire  _decoded_decoded_orMatrixOutputs_T_152 = |_decoded_decoded_T_57;
  wire  _decoded_decoded_orMatrixOutputs_T_153 = |_decoded_decoded_T_369;
  wire  _decoded_decoded_orMatrixOutputs_T_154 = |_decoded_decoded_T_245;
  wire  _decoded_decoded_orMatrixOutputs_T_155 = |_decoded_decoded_T_307;
  wire  _decoded_decoded_orMatrixOutputs_T_156 = |_decoded_decoded_T_183;
  wire  _decoded_decoded_orMatrixOutputs_T_157 = |_decoded_decoded_T_55;
  wire  _decoded_decoded_orMatrixOutputs_T_158 = |_decoded_decoded_T_367;
  wire  _decoded_decoded_orMatrixOutputs_T_159 = |_decoded_decoded_T_243;
  wire  _decoded_decoded_orMatrixOutputs_T_160 = |_decoded_decoded_T_305;
  wire  _decoded_decoded_orMatrixOutputs_T_161 = |_decoded_decoded_T_181;
  wire  _decoded_decoded_orMatrixOutputs_T_162 = |_decoded_decoded_T_53;
  wire  _decoded_decoded_orMatrixOutputs_T_163 = |_decoded_decoded_T_365;
  wire  _decoded_decoded_orMatrixOutputs_T_164 = |_decoded_decoded_T_241;
  wire  _decoded_decoded_orMatrixOutputs_T_165 = |_decoded_decoded_T_303;
  wire  _decoded_decoded_orMatrixOutputs_T_166 = |_decoded_decoded_T_179;
  wire  _decoded_decoded_orMatrixOutputs_T_167 = |_decoded_decoded_T_51;
  wire  _decoded_decoded_orMatrixOutputs_T_168 = |_decoded_decoded_T_363;
  wire  _decoded_decoded_orMatrixOutputs_T_169 = |_decoded_decoded_T_239;
  wire  _decoded_decoded_orMatrixOutputs_T_170 = |_decoded_decoded_T_301;
  wire  _decoded_decoded_orMatrixOutputs_T_171 = |_decoded_decoded_T_177;
  wire  _decoded_decoded_orMatrixOutputs_T_172 = |_decoded_decoded_T_49;
  wire  _decoded_decoded_orMatrixOutputs_T_173 = |_decoded_decoded_T_361;
  wire  _decoded_decoded_orMatrixOutputs_T_174 = |_decoded_decoded_T_237;
  wire  _decoded_decoded_orMatrixOutputs_T_175 = |_decoded_decoded_T_299;
  wire  _decoded_decoded_orMatrixOutputs_T_176 = |_decoded_decoded_T_175;
  wire  _decoded_decoded_orMatrixOutputs_T_177 = |_decoded_decoded_T_47;
  wire  _decoded_decoded_orMatrixOutputs_T_178 = |_decoded_decoded_T_359;
  wire  _decoded_decoded_orMatrixOutputs_T_179 = |_decoded_decoded_T_235;
  wire  _decoded_decoded_orMatrixOutputs_T_180 = |_decoded_decoded_T_297;
  wire  _decoded_decoded_orMatrixOutputs_T_181 = |_decoded_decoded_T_173;
  wire  _decoded_decoded_orMatrixOutputs_T_182 = |_decoded_decoded_T_45;
  wire  _decoded_decoded_orMatrixOutputs_T_183 = |_decoded_decoded_T_357;
  wire  _decoded_decoded_orMatrixOutputs_T_184 = |_decoded_decoded_T_233;
  wire  _decoded_decoded_orMatrixOutputs_T_185 = |_decoded_decoded_T_295;
  wire  _decoded_decoded_orMatrixOutputs_T_186 = |_decoded_decoded_T_171;
  wire  _decoded_decoded_orMatrixOutputs_T_187 = |_decoded_decoded_T_43;
  wire  _decoded_decoded_orMatrixOutputs_T_188 = |_decoded_decoded_T_169;
  wire  _decoded_decoded_orMatrixOutputs_T_189 = |_decoded_decoded_T_167;
  wire  _decoded_decoded_orMatrixOutputs_T_190 = |_decoded_decoded_T_41;
  wire  _decoded_decoded_orMatrixOutputs_T_191 = |_decoded_decoded_T_5;
  wire  _decoded_decoded_orMatrixOutputs_T_192 = |_decoded_decoded_T_3;
  wire  _decoded_decoded_orMatrixOutputs_T_193 = |_decoded_decoded_T_1;
  wire  _decoded_decoded_orMatrixOutputs_T_194 = |_decoded_decoded_T_163;
  wire  _decoded_decoded_orMatrixOutputs_T_195 = |_decoded_decoded_T_161;
  wire  _decoded_decoded_orMatrixOutputs_T_196 = |_decoded_decoded_T_159;
  wire  _decoded_decoded_orMatrixOutputs_T_197 = |_decoded_decoded_T_421;
  wire  _decoded_decoded_orMatrixOutputs_T_198 = |_decoded_decoded_T_105;
  wire  _decoded_decoded_orMatrixOutputs_T_199 = |_decoded_decoded_T_107;
  wire  _decoded_decoded_orMatrixOutputs_T_200 = |_decoded_decoded_T_103;
  wire  _decoded_decoded_orMatrixOutputs_T_201 = |_decoded_decoded_T_101;
  wire  _decoded_decoded_orMatrixOutputs_T_202 = |_decoded_decoded_T_35;
  wire  _decoded_decoded_orMatrixOutputs_T_203 = |_decoded_decoded_T_109;
  wire  _decoded_decoded_orMatrixOutputs_T_204 = |_decoded_decoded_T_37;
  wire  _decoded_decoded_orMatrixOutputs_T_205 = |_decoded_decoded_T_27;
  wire  _decoded_decoded_orMatrixOutputs_T_206 = |_decoded_decoded_T_29;
  wire  _decoded_decoded_orMatrixOutputs_T_207 = |_decoded_decoded_T_157;
  wire  _decoded_decoded_orMatrixOutputs_T_208 = |_decoded_decoded_T_155;
  wire  _decoded_decoded_orMatrixOutputs_T_209 = |_decoded_decoded_T_153;
  wire  _decoded_decoded_orMatrixOutputs_T_210 = |_decoded_decoded_T_151;
  wire [5:0] decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_5,
    _decoded_decoded_orMatrixOutputs_T_4,_decoded_decoded_orMatrixOutputs_T_3,_decoded_decoded_orMatrixOutputs_T_2,
    _decoded_decoded_orMatrixOutputs_T_1,_decoded_decoded_orMatrixOutputs_T};
  wire [12:0] decoded_decoded_orMatrixOutputs_lo_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_12,
    _decoded_decoded_orMatrixOutputs_T_11,_decoded_decoded_orMatrixOutputs_T_10,_decoded_decoded_orMatrixOutputs_T_9,
    _decoded_decoded_orMatrixOutputs_T_8,_decoded_decoded_orMatrixOutputs_T_7,_decoded_decoded_orMatrixOutputs_T_6,
    decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_18,
    _decoded_decoded_orMatrixOutputs_T_17,_decoded_decoded_orMatrixOutputs_T_16,_decoded_decoded_orMatrixOutputs_T_15,
    _decoded_decoded_orMatrixOutputs_T_14,_decoded_decoded_orMatrixOutputs_T_13};
  wire [25:0] decoded_decoded_orMatrixOutputs_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_25,
    _decoded_decoded_orMatrixOutputs_T_24,_decoded_decoded_orMatrixOutputs_T_23,_decoded_decoded_orMatrixOutputs_T_22,
    _decoded_decoded_orMatrixOutputs_T_21,_decoded_decoded_orMatrixOutputs_T_20,_decoded_decoded_orMatrixOutputs_T_19,
    decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo,decoded_decoded_orMatrixOutputs_lo_lo_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_31,
    _decoded_decoded_orMatrixOutputs_T_30,_decoded_decoded_orMatrixOutputs_T_29,_decoded_decoded_orMatrixOutputs_T_28,
    _decoded_decoded_orMatrixOutputs_T_27,_decoded_decoded_orMatrixOutputs_T_26};
  wire [12:0] decoded_decoded_orMatrixOutputs_lo_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_38,
    _decoded_decoded_orMatrixOutputs_T_37,_decoded_decoded_orMatrixOutputs_T_36,_decoded_decoded_orMatrixOutputs_T_35,
    _decoded_decoded_orMatrixOutputs_T_34,_decoded_decoded_orMatrixOutputs_T_33,_decoded_decoded_orMatrixOutputs_T_32,
    decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_44,
    _decoded_decoded_orMatrixOutputs_T_43,_decoded_decoded_orMatrixOutputs_T_42,_decoded_decoded_orMatrixOutputs_T_41,
    _decoded_decoded_orMatrixOutputs_T_40,_decoded_decoded_orMatrixOutputs_T_39};
  wire [51:0] decoded_decoded_orMatrixOutputs_lo_lo = {_decoded_decoded_orMatrixOutputs_T_51,
    _decoded_decoded_orMatrixOutputs_T_50,_decoded_decoded_orMatrixOutputs_T_49,_decoded_decoded_orMatrixOutputs_T_48,
    _decoded_decoded_orMatrixOutputs_T_47,_decoded_decoded_orMatrixOutputs_T_46,_decoded_decoded_orMatrixOutputs_T_45,
    decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo,decoded_decoded_orMatrixOutputs_lo_lo_hi_lo,
    decoded_decoded_orMatrixOutputs_lo_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_57,
    _decoded_decoded_orMatrixOutputs_T_56,_decoded_decoded_orMatrixOutputs_T_55,_decoded_decoded_orMatrixOutputs_T_54,
    _decoded_decoded_orMatrixOutputs_T_53,_decoded_decoded_orMatrixOutputs_T_52};
  wire [12:0] decoded_decoded_orMatrixOutputs_lo_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_64,
    _decoded_decoded_orMatrixOutputs_T_63,_decoded_decoded_orMatrixOutputs_T_62,_decoded_decoded_orMatrixOutputs_T_61,
    _decoded_decoded_orMatrixOutputs_T_60,_decoded_decoded_orMatrixOutputs_T_59,_decoded_decoded_orMatrixOutputs_T_58,
    decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_70,
    _decoded_decoded_orMatrixOutputs_T_69,_decoded_decoded_orMatrixOutputs_T_68,_decoded_decoded_orMatrixOutputs_T_67,
    _decoded_decoded_orMatrixOutputs_T_66,_decoded_decoded_orMatrixOutputs_T_65};
  wire [25:0] decoded_decoded_orMatrixOutputs_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_77,
    _decoded_decoded_orMatrixOutputs_T_76,_decoded_decoded_orMatrixOutputs_T_75,_decoded_decoded_orMatrixOutputs_T_74,
    _decoded_decoded_orMatrixOutputs_T_73,_decoded_decoded_orMatrixOutputs_T_72,_decoded_decoded_orMatrixOutputs_T_71,
    decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo,decoded_decoded_orMatrixOutputs_lo_hi_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_83,
    _decoded_decoded_orMatrixOutputs_T_82,_decoded_decoded_orMatrixOutputs_T_81,_decoded_decoded_orMatrixOutputs_T_80,
    _decoded_decoded_orMatrixOutputs_T_79,_decoded_decoded_orMatrixOutputs_T_78};
  wire [12:0] decoded_decoded_orMatrixOutputs_lo_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_90,
    _decoded_decoded_orMatrixOutputs_T_89,_decoded_decoded_orMatrixOutputs_T_88,_decoded_decoded_orMatrixOutputs_T_87,
    _decoded_decoded_orMatrixOutputs_T_86,_decoded_decoded_orMatrixOutputs_T_85,_decoded_decoded_orMatrixOutputs_T_84,
    decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo};
  wire [6:0] decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_97,
    _decoded_decoded_orMatrixOutputs_T_96,_decoded_decoded_orMatrixOutputs_T_95,_decoded_decoded_orMatrixOutputs_T_94,
    _decoded_decoded_orMatrixOutputs_T_93,_decoded_decoded_orMatrixOutputs_T_92,_decoded_decoded_orMatrixOutputs_T_91};
  wire [52:0] decoded_decoded_orMatrixOutputs_lo_hi = {_decoded_decoded_orMatrixOutputs_T_104,
    _decoded_decoded_orMatrixOutputs_T_103,_decoded_decoded_orMatrixOutputs_T_102,_decoded_decoded_orMatrixOutputs_T_101
    ,_decoded_decoded_orMatrixOutputs_T_100,_decoded_decoded_orMatrixOutputs_T_99,_decoded_decoded_orMatrixOutputs_T_98,
    decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo,decoded_decoded_orMatrixOutputs_lo_hi_hi_lo,
    decoded_decoded_orMatrixOutputs_lo_hi_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_110,
    _decoded_decoded_orMatrixOutputs_T_109,_decoded_decoded_orMatrixOutputs_T_108,_decoded_decoded_orMatrixOutputs_T_107
    ,_decoded_decoded_orMatrixOutputs_T_106,_decoded_decoded_orMatrixOutputs_T_105};
  wire [12:0] decoded_decoded_orMatrixOutputs_hi_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_117,
    _decoded_decoded_orMatrixOutputs_T_116,_decoded_decoded_orMatrixOutputs_T_115,_decoded_decoded_orMatrixOutputs_T_114
    ,_decoded_decoded_orMatrixOutputs_T_113,_decoded_decoded_orMatrixOutputs_T_112,
    _decoded_decoded_orMatrixOutputs_T_111,decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_123,
    _decoded_decoded_orMatrixOutputs_T_122,_decoded_decoded_orMatrixOutputs_T_121,_decoded_decoded_orMatrixOutputs_T_120
    ,_decoded_decoded_orMatrixOutputs_T_119,_decoded_decoded_orMatrixOutputs_T_118};
  wire [25:0] decoded_decoded_orMatrixOutputs_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_130,
    _decoded_decoded_orMatrixOutputs_T_129,_decoded_decoded_orMatrixOutputs_T_128,_decoded_decoded_orMatrixOutputs_T_127
    ,_decoded_decoded_orMatrixOutputs_T_126,_decoded_decoded_orMatrixOutputs_T_125,
    _decoded_decoded_orMatrixOutputs_T_124,decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo,
    decoded_decoded_orMatrixOutputs_hi_lo_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_136,
    _decoded_decoded_orMatrixOutputs_T_135,_decoded_decoded_orMatrixOutputs_T_134,_decoded_decoded_orMatrixOutputs_T_133
    ,_decoded_decoded_orMatrixOutputs_T_132,_decoded_decoded_orMatrixOutputs_T_131};
  wire [12:0] decoded_decoded_orMatrixOutputs_hi_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_143,
    _decoded_decoded_orMatrixOutputs_T_142,_decoded_decoded_orMatrixOutputs_T_141,_decoded_decoded_orMatrixOutputs_T_140
    ,_decoded_decoded_orMatrixOutputs_T_139,_decoded_decoded_orMatrixOutputs_T_138,
    _decoded_decoded_orMatrixOutputs_T_137,decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo};
  wire [6:0] decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_150,
    _decoded_decoded_orMatrixOutputs_T_149,_decoded_decoded_orMatrixOutputs_T_148,_decoded_decoded_orMatrixOutputs_T_147
    ,_decoded_decoded_orMatrixOutputs_T_146,_decoded_decoded_orMatrixOutputs_T_145,
    _decoded_decoded_orMatrixOutputs_T_144};
  wire [52:0] decoded_decoded_orMatrixOutputs_hi_lo = {_decoded_decoded_orMatrixOutputs_T_157,
    _decoded_decoded_orMatrixOutputs_T_156,_decoded_decoded_orMatrixOutputs_T_155,_decoded_decoded_orMatrixOutputs_T_154
    ,_decoded_decoded_orMatrixOutputs_T_153,_decoded_decoded_orMatrixOutputs_T_152,
    _decoded_decoded_orMatrixOutputs_T_151,decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo,
    decoded_decoded_orMatrixOutputs_hi_lo_hi_lo,decoded_decoded_orMatrixOutputs_hi_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_163,
    _decoded_decoded_orMatrixOutputs_T_162,_decoded_decoded_orMatrixOutputs_T_161,_decoded_decoded_orMatrixOutputs_T_160
    ,_decoded_decoded_orMatrixOutputs_T_159,_decoded_decoded_orMatrixOutputs_T_158};
  wire [12:0] decoded_decoded_orMatrixOutputs_hi_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_170,
    _decoded_decoded_orMatrixOutputs_T_169,_decoded_decoded_orMatrixOutputs_T_168,_decoded_decoded_orMatrixOutputs_T_167
    ,_decoded_decoded_orMatrixOutputs_T_166,_decoded_decoded_orMatrixOutputs_T_165,
    _decoded_decoded_orMatrixOutputs_T_164,decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_176,
    _decoded_decoded_orMatrixOutputs_T_175,_decoded_decoded_orMatrixOutputs_T_174,_decoded_decoded_orMatrixOutputs_T_173
    ,_decoded_decoded_orMatrixOutputs_T_172,_decoded_decoded_orMatrixOutputs_T_171};
  wire [25:0] decoded_decoded_orMatrixOutputs_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_183,
    _decoded_decoded_orMatrixOutputs_T_182,_decoded_decoded_orMatrixOutputs_T_181,_decoded_decoded_orMatrixOutputs_T_180
    ,_decoded_decoded_orMatrixOutputs_T_179,_decoded_decoded_orMatrixOutputs_T_178,
    _decoded_decoded_orMatrixOutputs_T_177,decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo,
    decoded_decoded_orMatrixOutputs_hi_hi_lo_lo};
  wire [5:0] decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_189,
    _decoded_decoded_orMatrixOutputs_T_188,_decoded_decoded_orMatrixOutputs_T_187,_decoded_decoded_orMatrixOutputs_T_186
    ,_decoded_decoded_orMatrixOutputs_T_185,_decoded_decoded_orMatrixOutputs_T_184};
  wire [12:0] decoded_decoded_orMatrixOutputs_hi_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_196,
    _decoded_decoded_orMatrixOutputs_T_195,_decoded_decoded_orMatrixOutputs_T_194,_decoded_decoded_orMatrixOutputs_T_193
    ,_decoded_decoded_orMatrixOutputs_T_192,_decoded_decoded_orMatrixOutputs_T_191,
    _decoded_decoded_orMatrixOutputs_T_190,decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo};
  wire [6:0] decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_203,
    _decoded_decoded_orMatrixOutputs_T_202,_decoded_decoded_orMatrixOutputs_T_201,_decoded_decoded_orMatrixOutputs_T_200
    ,_decoded_decoded_orMatrixOutputs_T_199,_decoded_decoded_orMatrixOutputs_T_198,
    _decoded_decoded_orMatrixOutputs_T_197};
  wire [52:0] decoded_decoded_orMatrixOutputs_hi_hi = {_decoded_decoded_orMatrixOutputs_T_210,
    _decoded_decoded_orMatrixOutputs_T_209,_decoded_decoded_orMatrixOutputs_T_208,_decoded_decoded_orMatrixOutputs_T_207
    ,_decoded_decoded_orMatrixOutputs_T_206,_decoded_decoded_orMatrixOutputs_T_205,
    _decoded_decoded_orMatrixOutputs_T_204,decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo,
    decoded_decoded_orMatrixOutputs_hi_hi_hi_lo,decoded_decoded_orMatrixOutputs_hi_hi_lo};
  wire [210:0] decoded_decoded_orMatrixOutputs = {decoded_decoded_orMatrixOutputs_hi_hi,
    decoded_decoded_orMatrixOutputs_hi_lo,decoded_decoded_orMatrixOutputs_lo_hi,decoded_decoded_orMatrixOutputs_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo = {decoded_decoded_orMatrixOutputs[5],
    decoded_decoded_orMatrixOutputs[4],decoded_decoded_orMatrixOutputs[3],decoded_decoded_orMatrixOutputs[2],
    decoded_decoded_orMatrixOutputs[1],decoded_decoded_orMatrixOutputs[0]};
  wire [12:0] decoded_decoded_invMatrixOutputs_lo_lo_lo_lo = {decoded_decoded_orMatrixOutputs[12],
    decoded_decoded_orMatrixOutputs[11],decoded_decoded_orMatrixOutputs[10],decoded_decoded_orMatrixOutputs[9],
    decoded_decoded_orMatrixOutputs[8],decoded_decoded_orMatrixOutputs[7],decoded_decoded_orMatrixOutputs[6],
    decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo = {decoded_decoded_orMatrixOutputs[18],
    decoded_decoded_orMatrixOutputs[17],decoded_decoded_orMatrixOutputs[16],decoded_decoded_orMatrixOutputs[15],
    decoded_decoded_orMatrixOutputs[14],decoded_decoded_orMatrixOutputs[13]};
  wire [25:0] decoded_decoded_invMatrixOutputs_lo_lo_lo = {decoded_decoded_orMatrixOutputs[25],
    decoded_decoded_orMatrixOutputs[24],decoded_decoded_orMatrixOutputs[23],decoded_decoded_orMatrixOutputs[22],
    decoded_decoded_orMatrixOutputs[21],decoded_decoded_orMatrixOutputs[20],decoded_decoded_orMatrixOutputs[19],
    decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo,decoded_decoded_invMatrixOutputs_lo_lo_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo = {decoded_decoded_orMatrixOutputs[31],
    decoded_decoded_orMatrixOutputs[30],decoded_decoded_orMatrixOutputs[29],decoded_decoded_orMatrixOutputs[28],
    decoded_decoded_orMatrixOutputs[27],decoded_decoded_orMatrixOutputs[26]};
  wire [12:0] decoded_decoded_invMatrixOutputs_lo_lo_hi_lo = {decoded_decoded_orMatrixOutputs[38],
    decoded_decoded_orMatrixOutputs[37],decoded_decoded_orMatrixOutputs[36],decoded_decoded_orMatrixOutputs[35],
    decoded_decoded_orMatrixOutputs[34],decoded_decoded_orMatrixOutputs[33],decoded_decoded_orMatrixOutputs[32],
    decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo = {decoded_decoded_orMatrixOutputs[44],
    decoded_decoded_orMatrixOutputs[43],decoded_decoded_orMatrixOutputs[42],decoded_decoded_orMatrixOutputs[41],
    decoded_decoded_orMatrixOutputs[40],decoded_decoded_orMatrixOutputs[39]};
  wire [51:0] decoded_decoded_invMatrixOutputs_lo_lo = {decoded_decoded_orMatrixOutputs[51],
    decoded_decoded_orMatrixOutputs[50],decoded_decoded_orMatrixOutputs[49],decoded_decoded_orMatrixOutputs[48],
    decoded_decoded_orMatrixOutputs[47],decoded_decoded_orMatrixOutputs[46],decoded_decoded_orMatrixOutputs[45],
    decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo,decoded_decoded_invMatrixOutputs_lo_lo_hi_lo,
    decoded_decoded_invMatrixOutputs_lo_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo = {decoded_decoded_orMatrixOutputs[57],
    decoded_decoded_orMatrixOutputs[56],decoded_decoded_orMatrixOutputs[55],decoded_decoded_orMatrixOutputs[54],
    decoded_decoded_orMatrixOutputs[53],decoded_decoded_orMatrixOutputs[52]};
  wire [12:0] decoded_decoded_invMatrixOutputs_lo_hi_lo_lo = {decoded_decoded_orMatrixOutputs[64],
    decoded_decoded_orMatrixOutputs[63],decoded_decoded_orMatrixOutputs[62],decoded_decoded_orMatrixOutputs[61],
    decoded_decoded_orMatrixOutputs[60],decoded_decoded_orMatrixOutputs[59],decoded_decoded_orMatrixOutputs[58],
    decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo = {decoded_decoded_orMatrixOutputs[70],
    decoded_decoded_orMatrixOutputs[69],decoded_decoded_orMatrixOutputs[68],decoded_decoded_orMatrixOutputs[67],
    decoded_decoded_orMatrixOutputs[66],decoded_decoded_orMatrixOutputs[65]};
  wire [25:0] decoded_decoded_invMatrixOutputs_lo_hi_lo = {decoded_decoded_orMatrixOutputs[77],
    decoded_decoded_orMatrixOutputs[76],decoded_decoded_orMatrixOutputs[75],decoded_decoded_orMatrixOutputs[74],
    decoded_decoded_orMatrixOutputs[73],decoded_decoded_orMatrixOutputs[72],decoded_decoded_orMatrixOutputs[71],
    decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo,decoded_decoded_invMatrixOutputs_lo_hi_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo = {decoded_decoded_orMatrixOutputs[83],
    decoded_decoded_orMatrixOutputs[82],decoded_decoded_orMatrixOutputs[81],decoded_decoded_orMatrixOutputs[80],
    decoded_decoded_orMatrixOutputs[79],decoded_decoded_orMatrixOutputs[78]};
  wire [12:0] decoded_decoded_invMatrixOutputs_lo_hi_hi_lo = {decoded_decoded_orMatrixOutputs[90],
    decoded_decoded_orMatrixOutputs[89],decoded_decoded_orMatrixOutputs[88],decoded_decoded_orMatrixOutputs[87],
    decoded_decoded_orMatrixOutputs[86],decoded_decoded_orMatrixOutputs[85],decoded_decoded_orMatrixOutputs[84],
    decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo};
  wire [6:0] decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo = {decoded_decoded_orMatrixOutputs[97],
    decoded_decoded_orMatrixOutputs[96],decoded_decoded_orMatrixOutputs[95],decoded_decoded_orMatrixOutputs[94],
    decoded_decoded_orMatrixOutputs[93],decoded_decoded_orMatrixOutputs[92],decoded_decoded_orMatrixOutputs[91]};
  wire [52:0] decoded_decoded_invMatrixOutputs_lo_hi = {decoded_decoded_orMatrixOutputs[104],
    decoded_decoded_orMatrixOutputs[103],decoded_decoded_orMatrixOutputs[102],decoded_decoded_orMatrixOutputs[101],
    decoded_decoded_orMatrixOutputs[100],decoded_decoded_orMatrixOutputs[99],decoded_decoded_orMatrixOutputs[98],
    decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo,decoded_decoded_invMatrixOutputs_lo_hi_hi_lo,
    decoded_decoded_invMatrixOutputs_lo_hi_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo = {decoded_decoded_orMatrixOutputs[110],
    decoded_decoded_orMatrixOutputs[109],decoded_decoded_orMatrixOutputs[108],decoded_decoded_orMatrixOutputs[107],
    decoded_decoded_orMatrixOutputs[106],decoded_decoded_orMatrixOutputs[105]};
  wire [12:0] decoded_decoded_invMatrixOutputs_hi_lo_lo_lo = {decoded_decoded_orMatrixOutputs[117],
    decoded_decoded_orMatrixOutputs[116],decoded_decoded_orMatrixOutputs[115],decoded_decoded_orMatrixOutputs[114],
    decoded_decoded_orMatrixOutputs[113],decoded_decoded_orMatrixOutputs[112],decoded_decoded_orMatrixOutputs[111],
    decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo = {decoded_decoded_orMatrixOutputs[123],
    decoded_decoded_orMatrixOutputs[122],decoded_decoded_orMatrixOutputs[121],decoded_decoded_orMatrixOutputs[120],
    decoded_decoded_orMatrixOutputs[119],decoded_decoded_orMatrixOutputs[118]};
  wire [25:0] decoded_decoded_invMatrixOutputs_hi_lo_lo = {decoded_decoded_orMatrixOutputs[130],
    decoded_decoded_orMatrixOutputs[129],decoded_decoded_orMatrixOutputs[128],decoded_decoded_orMatrixOutputs[127],
    decoded_decoded_orMatrixOutputs[126],decoded_decoded_orMatrixOutputs[125],decoded_decoded_orMatrixOutputs[124],
    decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo,decoded_decoded_invMatrixOutputs_hi_lo_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo = {decoded_decoded_orMatrixOutputs[136],
    decoded_decoded_orMatrixOutputs[135],decoded_decoded_orMatrixOutputs[134],decoded_decoded_orMatrixOutputs[133],
    decoded_decoded_orMatrixOutputs[132],decoded_decoded_orMatrixOutputs[131]};
  wire [12:0] decoded_decoded_invMatrixOutputs_hi_lo_hi_lo = {decoded_decoded_orMatrixOutputs[143],
    decoded_decoded_orMatrixOutputs[142],decoded_decoded_orMatrixOutputs[141],decoded_decoded_orMatrixOutputs[140],
    decoded_decoded_orMatrixOutputs[139],decoded_decoded_orMatrixOutputs[138],decoded_decoded_orMatrixOutputs[137],
    decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo};
  wire [6:0] decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo = {decoded_decoded_orMatrixOutputs[150],
    decoded_decoded_orMatrixOutputs[149],decoded_decoded_orMatrixOutputs[148],decoded_decoded_orMatrixOutputs[147],
    decoded_decoded_orMatrixOutputs[146],decoded_decoded_orMatrixOutputs[145],decoded_decoded_orMatrixOutputs[144]};
  wire [52:0] decoded_decoded_invMatrixOutputs_hi_lo = {decoded_decoded_orMatrixOutputs[157],
    decoded_decoded_orMatrixOutputs[156],decoded_decoded_orMatrixOutputs[155],decoded_decoded_orMatrixOutputs[154],
    decoded_decoded_orMatrixOutputs[153],decoded_decoded_orMatrixOutputs[152],decoded_decoded_orMatrixOutputs[151],
    decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo,decoded_decoded_invMatrixOutputs_hi_lo_hi_lo,
    decoded_decoded_invMatrixOutputs_hi_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo = {decoded_decoded_orMatrixOutputs[163],
    decoded_decoded_orMatrixOutputs[162],decoded_decoded_orMatrixOutputs[161],decoded_decoded_orMatrixOutputs[160],
    decoded_decoded_orMatrixOutputs[159],decoded_decoded_orMatrixOutputs[158]};
  wire [12:0] decoded_decoded_invMatrixOutputs_hi_hi_lo_lo = {decoded_decoded_orMatrixOutputs[170],
    decoded_decoded_orMatrixOutputs[169],decoded_decoded_orMatrixOutputs[168],decoded_decoded_orMatrixOutputs[167],
    decoded_decoded_orMatrixOutputs[166],decoded_decoded_orMatrixOutputs[165],decoded_decoded_orMatrixOutputs[164],
    decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo = {decoded_decoded_orMatrixOutputs[176],
    decoded_decoded_orMatrixOutputs[175],decoded_decoded_orMatrixOutputs[174],decoded_decoded_orMatrixOutputs[173],
    decoded_decoded_orMatrixOutputs[172],decoded_decoded_orMatrixOutputs[171]};
  wire [25:0] decoded_decoded_invMatrixOutputs_hi_hi_lo = {decoded_decoded_orMatrixOutputs[183],
    decoded_decoded_orMatrixOutputs[182],decoded_decoded_orMatrixOutputs[181],decoded_decoded_orMatrixOutputs[180],
    decoded_decoded_orMatrixOutputs[179],decoded_decoded_orMatrixOutputs[178],decoded_decoded_orMatrixOutputs[177],
    decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo,decoded_decoded_invMatrixOutputs_hi_hi_lo_lo};
  wire [5:0] decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo = {decoded_decoded_orMatrixOutputs[189],
    decoded_decoded_orMatrixOutputs[188],decoded_decoded_orMatrixOutputs[187],decoded_decoded_orMatrixOutputs[186],
    decoded_decoded_orMatrixOutputs[185],decoded_decoded_orMatrixOutputs[184]};
  wire [12:0] decoded_decoded_invMatrixOutputs_hi_hi_hi_lo = {decoded_decoded_orMatrixOutputs[196],
    decoded_decoded_orMatrixOutputs[195],decoded_decoded_orMatrixOutputs[194],decoded_decoded_orMatrixOutputs[193],
    decoded_decoded_orMatrixOutputs[192],decoded_decoded_orMatrixOutputs[191],decoded_decoded_orMatrixOutputs[190],
    decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo};
  wire [6:0] decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo = {decoded_decoded_orMatrixOutputs[203],
    decoded_decoded_orMatrixOutputs[202],decoded_decoded_orMatrixOutputs[201],decoded_decoded_orMatrixOutputs[200],
    decoded_decoded_orMatrixOutputs[199],decoded_decoded_orMatrixOutputs[198],decoded_decoded_orMatrixOutputs[197]};
  wire [52:0] decoded_decoded_invMatrixOutputs_hi_hi = {decoded_decoded_orMatrixOutputs[210],
    decoded_decoded_orMatrixOutputs[209],decoded_decoded_orMatrixOutputs[208],decoded_decoded_orMatrixOutputs[207],
    decoded_decoded_orMatrixOutputs[206],decoded_decoded_orMatrixOutputs[205],decoded_decoded_orMatrixOutputs[204],
    decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo,decoded_decoded_invMatrixOutputs_hi_hi_hi_lo,
    decoded_decoded_invMatrixOutputs_hi_hi_lo};
  wire [210:0] decoded_decoded_invMatrixOutputs = {decoded_decoded_invMatrixOutputs_hi_hi,
    decoded_decoded_invMatrixOutputs_hi_lo,decoded_decoded_invMatrixOutputs_lo_hi,decoded_decoded_invMatrixOutputs_lo_lo
    };
  wire  decoded_1 = decoded_decoded_invMatrixOutputs[209];
  wire  decoded_2 = decoded_decoded_invMatrixOutputs[208];
  wire  decoded_4 = decoded_decoded_invMatrixOutputs[206];
  wire  decoded_5 = decoded_decoded_invMatrixOutputs[205];
  wire  decoded_6 = decoded_decoded_invMatrixOutputs[204];
  wire  decoded_7 = decoded_decoded_invMatrixOutputs[203];
  wire  decoded_8 = decoded_decoded_invMatrixOutputs[202];
  wire  decoded_9 = decoded_decoded_invMatrixOutputs[201];
  wire  decoded_10 = decoded_decoded_invMatrixOutputs[200];
  wire  decoded_11 = decoded_decoded_invMatrixOutputs[199];
  wire  decoded_12 = decoded_decoded_invMatrixOutputs[198];
  wire  decoded_13 = decoded_decoded_invMatrixOutputs[197];
  wire  decoded_14 = decoded_decoded_invMatrixOutputs[196];
  wire  decoded_15 = decoded_decoded_invMatrixOutputs[195];
  wire  decoded_16 = decoded_decoded_invMatrixOutputs[194];
  wire  decoded_17 = decoded_decoded_invMatrixOutputs[193];
  wire  decoded_18 = decoded_decoded_invMatrixOutputs[192];
  wire  decoded_19 = decoded_decoded_invMatrixOutputs[191];
  wire  decoded_20 = decoded_decoded_invMatrixOutputs[190];
  wire  decoded_21 = decoded_decoded_invMatrixOutputs[189];
  wire  decoded_22 = decoded_decoded_invMatrixOutputs[188];
  wire  decoded_168 = decoded_decoded_invMatrixOutputs[42];
  wire  decoded_169 = decoded_decoded_invMatrixOutputs[41];
  wire  decoded_170 = decoded_decoded_invMatrixOutputs[40];
  wire  decoded_171 = decoded_decoded_invMatrixOutputs[39];
  wire  decoded_172 = decoded_decoded_invMatrixOutputs[38];
  wire  decoded_173 = decoded_decoded_invMatrixOutputs[37];
  wire  decoded_174 = decoded_decoded_invMatrixOutputs[36];
  wire  decoded_175 = decoded_decoded_invMatrixOutputs[35];
  wire  decoded_176 = decoded_decoded_invMatrixOutputs[34];
  wire  decoded_177 = decoded_decoded_invMatrixOutputs[33];
  wire  decoded_178 = decoded_decoded_invMatrixOutputs[32];
  wire  decoded_179 = decoded_decoded_invMatrixOutputs[31];
  wire  decoded_180 = decoded_decoded_invMatrixOutputs[30];
  wire  decoded_181 = decoded_decoded_invMatrixOutputs[29];
  wire  decoded_182 = decoded_decoded_invMatrixOutputs[28];
  wire  decoded_183 = decoded_decoded_invMatrixOutputs[27];
  wire  decoded_184 = decoded_decoded_invMatrixOutputs[26];
  wire  decoded_185 = decoded_decoded_invMatrixOutputs[25];
  wire  decoded_186 = decoded_decoded_invMatrixOutputs[24];
  wire  decoded_187 = decoded_decoded_invMatrixOutputs[23];
  wire  decoded_188 = decoded_decoded_invMatrixOutputs[22];
  wire  decoded_191 = decoded_decoded_invMatrixOutputs[19];
  wire  decoded_192 = decoded_decoded_invMatrixOutputs[18];
  wire  decoded_193 = decoded_decoded_invMatrixOutputs[17];
  wire  decoded_194 = decoded_decoded_invMatrixOutputs[16];
  wire  decoded_195 = decoded_decoded_invMatrixOutputs[15];
  wire  decoded_196 = decoded_decoded_invMatrixOutputs[14];
  wire  decoded_197 = decoded_decoded_invMatrixOutputs[13];
  wire  decoded_198 = decoded_decoded_invMatrixOutputs[12];
  wire  decoded_207 = decoded_decoded_invMatrixOutputs[3];
  wire  decoded_208 = decoded_decoded_invMatrixOutputs[2];
  wire  decoded_210 = decoded_decoded_invMatrixOutputs[0];
  wire [31:0] _wdata_T_1 = io_rw_cmd[1] ? io_rw_rdata : 32'h0;
  wire [31:0] _wdata_T_2 = _wdata_T_1 | io_rw_wdata;
  wire [31:0] _wdata_T_5 = &io_rw_cmd[1:0] ? io_rw_wdata : 32'h0;
  wire [31:0] _wdata_T_6 = ~_wdata_T_5;
  wire [31:0] wdata = _wdata_T_2 & _wdata_T_6;
  wire  insn_cease = system_insn & decoded_invMatrixOutputs[5];
  wire  insn_wfi = system_insn & decoded_invMatrixOutputs[4];
  wire [11:0] addr_1 = io_decode_0_inst[31:20];
  wire [31:0] decoded_invInputs_1 = ~io_decode_0_inst;
  wire  decoded_andMatrixInput_0_7 = decoded_invInputs_1[20];
  wire  decoded_andMatrixInput_1_7 = decoded_invInputs_1[21];
  wire  decoded_andMatrixInput_2_6 = decoded_invInputs_1[22];
  wire  decoded_andMatrixInput_3_6 = decoded_invInputs_1[23];
  wire  decoded_andMatrixInput_4_6 = decoded_invInputs_1[24];
  wire  decoded_andMatrixInput_5_6 = decoded_invInputs_1[25];
  wire  decoded_andMatrixInput_6_6 = decoded_invInputs_1[26];
  wire  decoded_andMatrixInput_7_6 = decoded_invInputs_1[27];
  wire  decoded_andMatrixInput_8_6 = decoded_invInputs_1[28];
  wire  decoded_andMatrixInput_9_6 = decoded_invInputs_1[29];
  wire  decoded_andMatrixInput_10_3 = decoded_invInputs_1[30];
  wire  decoded_andMatrixInput_11_3 = decoded_invInputs_1[31];
  wire [5:0] decoded_lo_6 = {decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,decoded_andMatrixInput_8_6,
    decoded_andMatrixInput_9_6,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3};
  wire [11:0] _decoded_T_14 = {decoded_andMatrixInput_0_7,decoded_andMatrixInput_1_7,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,decoded_andMatrixInput_5_6,decoded_lo_6};
  wire  _decoded_T_15 = &_decoded_T_14;
  wire  decoded_andMatrixInput_0_8 = io_decode_0_inst[20];
  wire [11:0] _decoded_T_16 = {decoded_andMatrixInput_0_8,decoded_andMatrixInput_1_7,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,decoded_andMatrixInput_5_6,decoded_lo_6};
  wire  _decoded_T_17 = &_decoded_T_16;
  wire  decoded_andMatrixInput_0_9 = io_decode_0_inst[0];
  wire  decoded_andMatrixInput_7_8 = io_decode_0_inst[28];
  wire [9:0] _decoded_T_18 = {decoded_andMatrixInput_0_9,decoded_andMatrixInput_2_6,decoded_andMatrixInput_3_6,
    decoded_andMatrixInput_4_6,decoded_andMatrixInput_5_6,decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,
    decoded_andMatrixInput_7_8,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3};
  wire  _decoded_T_19 = &_decoded_T_18;
  wire  decoded_andMatrixInput_0_10 = io_decode_0_inst[22];
  wire [9:0] _decoded_T_20 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,
    decoded_andMatrixInput_5_6,decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,decoded_andMatrixInput_7_8,
    decoded_andMatrixInput_9_6,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3};
  wire  _decoded_T_21 = &_decoded_T_20;
  wire  decoded_andMatrixInput_1_11 = io_decode_0_inst[1];
  wire  decoded_andMatrixInput_2_10 = decoded_invInputs_1[2];
  wire  decoded_andMatrixInput_3_10 = decoded_invInputs_1[3];
  wire  decoded_andMatrixInput_4_10 = io_decode_0_inst[4];
  wire  decoded_andMatrixInput_5_10 = io_decode_0_inst[5];
  wire  decoded_andMatrixInput_6_10 = io_decode_0_inst[6];
  wire  decoded_andMatrixInput_7_10 = decoded_invInputs_1[7];
  wire  decoded_andMatrixInput_8_10 = decoded_invInputs_1[8];
  wire  decoded_andMatrixInput_9_10 = decoded_invInputs_1[9];
  wire  decoded_andMatrixInput_10_5 = io_decode_0_inst[25];
  wire [7:0] decoded_lo_10 = {decoded_andMatrixInput_9_10,decoded_andMatrixInput_10_5,decoded_andMatrixInput_6_6,
    decoded_andMatrixInput_7_6,decoded_andMatrixInput_7_8,decoded_andMatrixInput_9_6,decoded_andMatrixInput_10_3,
    decoded_andMatrixInput_11_3};
  wire [16:0] _decoded_T_22 = {decoded_andMatrixInput_0_9,decoded_andMatrixInput_1_11,decoded_andMatrixInput_2_10,
    decoded_andMatrixInput_3_10,decoded_andMatrixInput_4_10,decoded_andMatrixInput_5_10,decoded_andMatrixInput_6_10,
    decoded_andMatrixInput_7_10,decoded_andMatrixInput_8_10,decoded_lo_10};
  wire  _decoded_T_23 = &_decoded_T_22;
  wire  decoded_andMatrixInput_7_11 = io_decode_0_inst[29];
  wire [9:0] _decoded_T_24 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,
    decoded_andMatrixInput_5_6,decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,decoded_andMatrixInput_7_8,
    decoded_andMatrixInput_7_11,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3};
  wire  _decoded_T_25 = &_decoded_T_24;
  wire  decoded_andMatrixInput_0_13 = io_decode_0_inst[30];
  wire [1:0] _decoded_T_26 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_11_3};
  wire  _decoded_T_27 = &_decoded_T_26;
  wire  _decoded_orMatrixOutputs_T_7 = |_decoded_T_23;
  wire  _decoded_orMatrixOutputs_T_8 = |_decoded_T_21;
  wire  _decoded_orMatrixOutputs_T_9 = |_decoded_T_25;
  wire [1:0] _decoded_orMatrixOutputs_T_10 = {_decoded_T_19,_decoded_T_27};
  wire  _decoded_orMatrixOutputs_T_11 = |_decoded_orMatrixOutputs_T_10;
  wire  _decoded_orMatrixOutputs_T_12 = |_decoded_T_17;
  wire  _decoded_orMatrixOutputs_T_13 = |_decoded_T_15;
  wire [8:0] decoded_orMatrixOutputs_1 = {_decoded_orMatrixOutputs_T_13,_decoded_orMatrixOutputs_T_12,
    _decoded_orMatrixOutputs_T_11,_decoded_orMatrixOutputs_T_9,_decoded_orMatrixOutputs_T_8,_decoded_orMatrixOutputs_T_7
    ,1'h0,2'h0};
  wire [8:0] decoded_invMatrixOutputs_1 = {decoded_orMatrixOutputs_1[8],decoded_orMatrixOutputs_1[7],
    decoded_orMatrixOutputs_1[6],decoded_orMatrixOutputs_1[5],decoded_orMatrixOutputs_1[4],decoded_orMatrixOutputs_1[3],
    decoded_orMatrixOutputs_1[2],decoded_orMatrixOutputs_1[1],decoded_orMatrixOutputs_1[0]};
  wire  is_ret = decoded_invMatrixOutputs_1[6];
  wire  is_wfi = decoded_invMatrixOutputs_1[4];
  wire  is_sfence = decoded_invMatrixOutputs_1[3];
  wire  is_hfence_gvma = decoded_invMatrixOutputs_1[1];
  wire  is_hlsv = decoded_invMatrixOutputs_1[0];
  wire  _is_counter_T_2 = addr_1 >= 12'hc00 & addr_1 < 12'hc20;
  wire  _is_counter_T_5 = addr_1 >= 12'hc80 & addr_1 < 12'hca0;
  wire  is_counter = _is_counter_T_2 | _is_counter_T_5;
  wire  _allow_wfi_T = reg_mstatus_prv > 2'h1;
  wire  allow_wfi = reg_mstatus_prv > 2'h1 | ~reg_mstatus_tw;
  wire  allow_sfence_vma = _allow_wfi_T | ~reg_mstatus_tvm;
  wire  _allow_hfence_vvma_T_1 = reg_mstatus_prv >= 2'h1;
  wire  allow_sret = _allow_wfi_T | ~reg_mstatus_tsr;
  wire [4:0] counter_addr = addr_1[4:0];
  wire [31:0] _allow_counter_T_1 = read_mcounteren >> counter_addr;
  wire [31:0] _allow_counter_T_6 = read_scounteren >> counter_addr;
  wire  _allow_counter_T_8 = _allow_hfence_vvma_T_1 | _allow_counter_T_6[0];
  wire  allow_counter = (_allow_wfi_T | _allow_counter_T_1[0]) & _allow_counter_T_8;
  wire [11:0] io_decode_0_fp_csr_invInputs = ~addr_1;
  wire  io_decode_0_fp_csr_andMatrixInput_0 = io_decode_0_fp_csr_invInputs[8];
  wire  io_decode_0_fp_csr_andMatrixInput_1 = io_decode_0_fp_csr_invInputs[9];
  wire  io_decode_0_fp_csr_andMatrixInput_2 = io_decode_0_fp_csr_invInputs[10];
  wire  io_decode_0_fp_csr_andMatrixInput_3 = io_decode_0_fp_csr_invInputs[11];
  wire [3:0] _io_decode_0_fp_csr_T = {io_decode_0_fp_csr_andMatrixInput_0,io_decode_0_fp_csr_andMatrixInput_1,
    io_decode_0_fp_csr_andMatrixInput_2,io_decode_0_fp_csr_andMatrixInput_3};
  wire  _io_decode_0_fp_csr_T_1 = &_io_decode_0_fp_csr_T;
  wire  csr_addr_legal = reg_mstatus_prv >= addr_1[9:8];
  wire  _csr_exists_T_15 = addr_1 == 12'h7b1;
  wire  _csr_exists_T_181 = addr_1 == 12'h180;
  wire  _csr_exists_T_225 = addr_1 == 12'h7a0 | addr_1 == 12'h7a1 | addr_1 == 12'h7a2 | addr_1 == 12'h7a3 | addr_1 == 12'h301
     | addr_1 == 12'h300 | addr_1 == 12'h305 | addr_1 == 12'h344 | addr_1 == 12'h304 | addr_1 == 12'h340 | addr_1 == 12'h341
     | addr_1 == 12'h343 | addr_1 == 12'h342 | addr_1 == 12'hf14 | addr_1 == 12'h7b0 | _csr_exists_T_15;
  wire  _csr_exists_T_240 = _csr_exists_T_225 | addr_1 == 12'h7b2 | addr_1 == 12'h1 | addr_1 == 12'h2 | addr_1 == 12'h3
     | addr_1 == 12'h320 | addr_1 == 12'hb00 | addr_1 == 12'hb02 | addr_1 == 12'h323 | addr_1 == 12'hb03 | addr_1 == 12'hc03
     | addr_1 == 12'hb83 | addr_1 == 12'hc83 | addr_1 == 12'h324 | addr_1 == 12'hb04 | addr_1 == 12'hc04;
  wire  _csr_exists_T_255 = _csr_exists_T_240 | addr_1 == 12'hb84 | addr_1 == 12'hc84 | addr_1 == 12'h325 | addr_1 == 12'hb05
     | addr_1 == 12'hc05 | addr_1 == 12'hb85 | addr_1 == 12'hc85 | addr_1 == 12'h326 | addr_1 == 12'hb06 | addr_1 == 12'hc06
     | addr_1 == 12'hb86 | addr_1 == 12'hc86 | addr_1 == 12'h327 | addr_1 == 12'hb07 | addr_1 == 12'hc07;
  wire  _csr_exists_T_270 = _csr_exists_T_255 | addr_1 == 12'hb87 | addr_1 == 12'hc87 | addr_1 == 12'h328 | addr_1 == 12'hb08
     | addr_1 == 12'hc08 | addr_1 == 12'hb88 | addr_1 == 12'hc88 | addr_1 == 12'h329 | addr_1 == 12'hb09 | addr_1 == 12'hc09
     | addr_1 == 12'hb89 | addr_1 == 12'hc89 | addr_1 == 12'h32a | addr_1 == 12'hb0a | addr_1 == 12'hc0a;
  wire  _csr_exists_T_285 = _csr_exists_T_270 | addr_1 == 12'hb8a | addr_1 == 12'hc8a | addr_1 == 12'h32b | addr_1 == 12'hb0b
     | addr_1 == 12'hc0b | addr_1 == 12'hb8b | addr_1 == 12'hc8b | addr_1 == 12'h32c | addr_1 == 12'hb0c | addr_1 == 12'hc0c
     | addr_1 == 12'hb8c | addr_1 == 12'hc8c | addr_1 == 12'h32d | addr_1 == 12'hb0d | addr_1 == 12'hc0d;
  wire  _csr_exists_T_300 = _csr_exists_T_285 | addr_1 == 12'hb8d | addr_1 == 12'hc8d | addr_1 == 12'h32e | addr_1 == 12'hb0e
     | addr_1 == 12'hc0e | addr_1 == 12'hb8e | addr_1 == 12'hc8e | addr_1 == 12'h32f | addr_1 == 12'hb0f | addr_1 == 12'hc0f
     | addr_1 == 12'hb8f | addr_1 == 12'hc8f | addr_1 == 12'h330 | addr_1 == 12'hb10 | addr_1 == 12'hc10;
  wire  _csr_exists_T_315 = _csr_exists_T_300 | addr_1 == 12'hb90 | addr_1 == 12'hc90 | addr_1 == 12'h331 | addr_1 == 12'hb11
     | addr_1 == 12'hc11 | addr_1 == 12'hb91 | addr_1 == 12'hc91 | addr_1 == 12'h332 | addr_1 == 12'hb12 | addr_1 == 12'hc12
     | addr_1 == 12'hb92 | addr_1 == 12'hc92 | addr_1 == 12'h333 | addr_1 == 12'hb13 | addr_1 == 12'hc13;
  wire  _csr_exists_T_330 = _csr_exists_T_315 | addr_1 == 12'hb93 | addr_1 == 12'hc93 | addr_1 == 12'h334 | addr_1 == 12'hb14
     | addr_1 == 12'hc14 | addr_1 == 12'hb94 | addr_1 == 12'hc94 | addr_1 == 12'h335 | addr_1 == 12'hb15 | addr_1 == 12'hc15
     | addr_1 == 12'hb95 | addr_1 == 12'hc95 | addr_1 == 12'h336 | addr_1 == 12'hb16 | addr_1 == 12'hc16;
  wire  _csr_exists_T_345 = _csr_exists_T_330 | addr_1 == 12'hb96 | addr_1 == 12'hc96 | addr_1 == 12'h337 | addr_1 == 12'hb17
     | addr_1 == 12'hc17 | addr_1 == 12'hb97 | addr_1 == 12'hc97 | addr_1 == 12'h338 | addr_1 == 12'hb18 | addr_1 == 12'hc18
     | addr_1 == 12'hb98 | addr_1 == 12'hc98 | addr_1 == 12'h339 | addr_1 == 12'hb19 | addr_1 == 12'hc19;
  wire  _csr_exists_T_360 = _csr_exists_T_345 | addr_1 == 12'hb99 | addr_1 == 12'hc99 | addr_1 == 12'h33a | addr_1 == 12'hb1a
     | addr_1 == 12'hc1a | addr_1 == 12'hb9a | addr_1 == 12'hc9a | addr_1 == 12'h33b | addr_1 == 12'hb1b | addr_1 == 12'hc1b
     | addr_1 == 12'hb9b | addr_1 == 12'hc9b | addr_1 == 12'h33c | addr_1 == 12'hb1c | addr_1 == 12'hc1c;
  wire  _csr_exists_T_375 = _csr_exists_T_360 | addr_1 == 12'hb9c | addr_1 == 12'hc9c | addr_1 == 12'h33d | addr_1 == 12'hb1d
     | addr_1 == 12'hc1d | addr_1 == 12'hb9d | addr_1 == 12'hc9d | addr_1 == 12'h33e | addr_1 == 12'hb1e | addr_1 == 12'hc1e
     | addr_1 == 12'hb9e | addr_1 == 12'hc9e | addr_1 == 12'h33f | addr_1 == 12'hb1f | addr_1 == 12'hc1f;
  wire  _csr_exists_T_390 = _csr_exists_T_375 | addr_1 == 12'hb9f | addr_1 == 12'hc9f | addr_1 == 12'h306 | addr_1 == 12'hc00
     | addr_1 == 12'hc02 | addr_1 == 12'hb80 | addr_1 == 12'hb82 | addr_1 == 12'hc80 | addr_1 == 12'hc82 | addr_1 == 12'h100
     | addr_1 == 12'h144 | addr_1 == 12'h104 | addr_1 == 12'h140 | addr_1 == 12'h142 | addr_1 == 12'h143;
  wire  _csr_exists_T_405 = _csr_exists_T_390 | addr_1 == 12'h180 | addr_1 == 12'h141 | addr_1 == 12'h105 | addr_1 == 12'h106
     | addr_1 == 12'h303 | addr_1 == 12'h302 | addr_1 == 12'h3a0 | addr_1 == 12'h3a1 | addr_1 == 12'h3a2 | addr_1 == 12'h3a3
     | addr_1 == 12'h3b0 | addr_1 == 12'h3b1 | addr_1 == 12'h3b2 | addr_1 == 12'h3b3 | addr_1 == 12'h3b4;
  wire  csr_exists = _csr_exists_T_405 | addr_1 == 12'h3b5 | addr_1 == 12'h3b6 | addr_1 == 12'h3b7 | addr_1 == 12'h3b8
     | addr_1 == 12'h3b9 | addr_1 == 12'h3ba | addr_1 == 12'h3bb | addr_1 == 12'h3bc | addr_1 == 12'h3bd | addr_1 == 12'h3be
     | addr_1 == 12'h3bf | addr_1 == 12'h7c1 | addr_1 == 12'hf12 | addr_1 == 12'hf11 | addr_1 == 12'hf13;
  wire  _io_decode_0_read_illegal_T = ~csr_addr_legal;
  wire  _io_decode_0_read_illegal_T_1 = ~csr_exists;
  wire  _io_decode_0_read_illegal_T_2 = ~csr_addr_legal | _io_decode_0_read_illegal_T_1;
  wire  _io_decode_0_read_illegal_T_6 = ~allow_sfence_vma;
  wire  _io_decode_0_read_illegal_T_7 = (_csr_exists_T_181 | addr_1 == 12'h680) & ~allow_sfence_vma;
  wire  _io_decode_0_read_illegal_T_8 = _io_decode_0_read_illegal_T_2 | _io_decode_0_read_illegal_T_7;
  wire  _io_decode_0_read_illegal_T_10 = is_counter & ~allow_counter;
  wire  _io_decode_0_read_illegal_T_11 = _io_decode_0_read_illegal_T_8 | _io_decode_0_read_illegal_T_10;
  wire  io_decode_0_read_illegal_andMatrixInput_0 = addr_1[4];
  wire  io_decode_0_read_illegal_andMatrixInput_1 = addr_1[5];
  wire  io_decode_0_read_illegal_andMatrixInput_2 = io_decode_0_fp_csr_invInputs[6];
  wire  io_decode_0_read_illegal_andMatrixInput_3 = addr_1[7];
  wire  io_decode_0_read_illegal_andMatrixInput_4 = addr_1[8];
  wire  io_decode_0_read_illegal_andMatrixInput_5 = addr_1[9];
  wire  io_decode_0_read_illegal_andMatrixInput_6 = addr_1[10];
  wire [7:0] _io_decode_0_read_illegal_T_12 = {io_decode_0_read_illegal_andMatrixInput_0,
    io_decode_0_read_illegal_andMatrixInput_1,io_decode_0_read_illegal_andMatrixInput_2,
    io_decode_0_read_illegal_andMatrixInput_3,io_decode_0_read_illegal_andMatrixInput_4,
    io_decode_0_read_illegal_andMatrixInput_5,io_decode_0_read_illegal_andMatrixInput_6,
    io_decode_0_fp_csr_andMatrixInput_3};
  wire  _io_decode_0_read_illegal_T_13 = &_io_decode_0_read_illegal_T_12;
  wire  io_decode_0_read_illegal_orMatrixOutputs = |_io_decode_0_read_illegal_T_13;
  wire  _io_decode_0_read_illegal_T_16 = io_decode_0_read_illegal_orMatrixOutputs & _T_397;
  wire  _io_decode_0_read_illegal_T_17 = _io_decode_0_read_illegal_T_11 | _io_decode_0_read_illegal_T_16;
  wire  _io_decode_0_read_illegal_T_21 = io_decode_0_fp_csr & io_decode_0_fp_illegal;
  wire [11:0] io_decode_0_write_flush_addr_m = addr_1 | 12'h300;
  wire  _io_decode_0_system_illegal_T_4 = is_wfi & ~allow_wfi;
  wire  _io_decode_0_system_illegal_T_5 = _io_decode_0_read_illegal_T & ~is_hlsv | _io_decode_0_system_illegal_T_4;
  wire  _io_decode_0_system_illegal_T_7 = is_ret & ~allow_sret;
  wire  _io_decode_0_system_illegal_T_8 = _io_decode_0_system_illegal_T_5 | _io_decode_0_system_illegal_T_7;
  wire  _io_decode_0_system_illegal_T_14 = is_ret & io_decode_0_read_illegal_andMatrixInput_6 &
    io_decode_0_read_illegal_andMatrixInput_3 & _T_397;
  wire  _io_decode_0_system_illegal_T_15 = _io_decode_0_system_illegal_T_8 | _io_decode_0_system_illegal_T_14;
  wire  _io_decode_0_system_illegal_T_18 = (is_sfence | is_hfence_gvma) & _io_decode_0_read_illegal_T_6;
  wire [11:0] _debugTVec_T = insn_break ? 12'h800 : 12'h808;
  wire [11:0] debugTVec = reg_debug ? _debugTVec_T : 12'h800;
  wire [31:0] notDebugTVec_base = delegate ? read_stvec : read_mtvec;
  wire [6:0] notDebugTVec_interruptOffset = {cause[4:0], 2'h0};
  wire [31:0] notDebugTVec_interruptVec = {notDebugTVec_base[31:7],notDebugTVec_interruptOffset};
  wire  notDebugTVec_doVector = notDebugTVec_base[0] & cause[31] & cause_lsbs[7:5] == 3'h0;
  wire [31:0] _notDebugTVec_T_1 = {notDebugTVec_base[31:2], 2'h0};
  wire [31:0] notDebugTVec = notDebugTVec_doVector ? notDebugTVec_interruptVec : _notDebugTVec_T_1;
  wire [31:0] tvec = trapToDebug ? {{20'd0}, debugTVec} : notDebugTVec;
  wire [1:0] _T_365 = insn_ret + insn_call;
  wire [1:0] _T_367 = insn_break + io_exception;
  wire [2:0] _T_369 = _T_365 + _T_367;
  wire  _T_373 = ~reset;
  wire  _GEN_46 = insn_wfi & _io_interrupt_T & _T_397 | reg_wfi;
  wire  _GEN_48 = io_retire | exception | reg_singleStepped;
  wire [31:0] _epc_T = ~io_pc;
  wire [31:0] _epc_T_1 = _epc_T | 32'h1;
  wire [31:0] epc = ~_epc_T_1;
  wire [1:0] _reg_dcsr_cause_T = causeIsDebugTrigger ? 2'h2 : 2'h1;
  wire [1:0] _reg_dcsr_cause_T_1 = causeIsDebugInt ? 2'h3 : _reg_dcsr_cause_T;
  wire [2:0] _reg_dcsr_cause_T_2 = reg_singleStepped ? 3'h4 : {{1'd0}, _reg_dcsr_cause_T_1};
  wire  _GEN_51 = ~reg_debug | reg_debug;
  wire [31:0] _GEN_52 = ~reg_debug ? epc : reg_dpc;
  wire [1:0] _GEN_54 = ~reg_debug ? reg_mstatus_prv : reg_dcsr_prv;
  wire [31:0] _GEN_68 = delegate ? epc : reg_sepc;
  wire [31:0] _GEN_69 = delegate ? cause : reg_scause;
  wire [31:0] _GEN_70 = delegate ? io_tval : reg_stval;
  wire  _GEN_72 = delegate ? reg_mstatus_sie : reg_mstatus_spie;
  wire [1:0] _GEN_73 = delegate ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp};
  wire  _GEN_74 = delegate ? 1'h0 : reg_mstatus_sie;
  wire [31:0] _GEN_78 = delegate ? reg_mepc : epc;
  wire [31:0] _GEN_79 = delegate ? reg_mcause : cause;
  wire [31:0] _GEN_80 = delegate ? reg_mtval : io_tval;
  wire  _GEN_82 = delegate ? reg_mstatus_mpie : reg_mstatus_mie;
  wire [1:0] _GEN_83 = delegate ? reg_mstatus_mpp : reg_mstatus_prv;
  wire  _GEN_84 = delegate & reg_mstatus_mie;
  wire  _GEN_145 = trapToDebug ? _GEN_51 : reg_debug;
  wire [31:0] _GEN_146 = trapToDebug ? _GEN_52 : reg_dpc;
  wire [1:0] _GEN_148 = trapToDebug ? _GEN_54 : reg_dcsr_prv;
  wire [31:0] _GEN_165 = trapToDebug ? reg_sepc : _GEN_68;
  wire [31:0] _GEN_166 = trapToDebug ? reg_scause : _GEN_69;
  wire [31:0] _GEN_167 = trapToDebug ? reg_stval : _GEN_70;
  wire  _GEN_169 = trapToDebug ? reg_mstatus_spie : _GEN_72;
  wire [1:0] _GEN_170 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_73;
  wire  _GEN_171 = trapToDebug ? reg_mstatus_sie : _GEN_74;
  wire [31:0] _GEN_174 = trapToDebug ? reg_mepc : _GEN_78;
  wire [31:0] _GEN_175 = trapToDebug ? reg_mcause : _GEN_79;
  wire [31:0] _GEN_176 = trapToDebug ? reg_mtval : _GEN_80;
  wire  _GEN_178 = trapToDebug ? reg_mstatus_mpie : _GEN_82;
  wire [1:0] _GEN_179 = trapToDebug ? reg_mstatus_mpp : _GEN_83;
  wire  _GEN_180 = trapToDebug ? reg_mstatus_mie : _GEN_84;
  wire  _GEN_182 = exception ? _GEN_145 : reg_debug;
  wire [31:0] _GEN_183 = exception ? _GEN_146 : reg_dpc;
  wire [1:0] _GEN_185 = exception ? _GEN_148 : reg_dcsr_prv;
  wire [31:0] _GEN_202 = exception ? _GEN_165 : reg_sepc;
  wire [31:0] _GEN_203 = exception ? _GEN_166 : reg_scause;
  wire [31:0] _GEN_204 = exception ? _GEN_167 : reg_stval;
  wire  _GEN_206 = exception ? _GEN_169 : reg_mstatus_spie;
  wire [1:0] _GEN_207 = exception ? _GEN_170 : {{1'd0}, reg_mstatus_spp};
  wire  _GEN_208 = exception ? _GEN_171 : reg_mstatus_sie;
  wire [31:0] _GEN_211 = exception ? _GEN_174 : reg_mepc;
  wire [31:0] _GEN_212 = exception ? _GEN_175 : reg_mcause;
  wire [31:0] _GEN_213 = exception ? _GEN_176 : reg_mtval;
  wire  _GEN_215 = exception ? _GEN_178 : reg_mstatus_mpie;
  wire [1:0] _GEN_216 = exception ? _GEN_179 : reg_mstatus_mpp;
  wire  _GEN_217 = exception ? _GEN_180 : reg_mstatus_mie;
  wire [31:0] _GEN_239 = io_rw_addr[10] & io_rw_addr[7] ? _T_28 : _T_22;
  wire  _GEN_241 = io_rw_addr[10] & io_rw_addr[7] ? _GEN_217 : reg_mstatus_mpie;
  wire  _GEN_242 = io_rw_addr[10] & io_rw_addr[7] ? _GEN_215 : 1'h1;
  wire [1:0] _GEN_243 = io_rw_addr[10] & io_rw_addr[7] ? _GEN_216 : 2'h0;
  wire  _GEN_245 = ~io_rw_addr[9] ? reg_mstatus_spie : _GEN_208;
  wire  _GEN_246 = ~io_rw_addr[9] | _GEN_206;
  wire [1:0] _GEN_247 = ~io_rw_addr[9] ? 2'h0 : _GEN_207;
  wire [31:0] _GEN_250 = ~io_rw_addr[9] ? _T_98 : _GEN_239;
  wire  _GEN_257 = ~io_rw_addr[9] ? _GEN_217 : _GEN_241;
  wire  _GEN_258 = ~io_rw_addr[9] ? _GEN_215 : _GEN_242;
  wire [1:0] _GEN_259 = ~io_rw_addr[9] ? _GEN_216 : _GEN_243;
  wire  _GEN_261 = ret_prv <= 2'h1 ? 1'h0 : reg_mstatus_mprv;
  wire  _GEN_262 = insn_ret ? _GEN_245 : _GEN_208;
  wire  _GEN_263 = insn_ret ? _GEN_246 : _GEN_206;
  wire [1:0] _GEN_264 = insn_ret ? _GEN_247 : _GEN_207;
  wire  _GEN_273 = insn_ret ? _GEN_257 : _GEN_217;
  wire  _GEN_274 = insn_ret ? _GEN_258 : _GEN_215;
  wire [1:0] _GEN_275 = insn_ret ? _GEN_259 : _GEN_216;
  wire  _GEN_278 = insn_ret ? _GEN_261 : reg_mstatus_mprv;
  reg  io_status_cease_r;
  wire  _GEN_279 = insn_cease | io_status_cease_r;
  wire [31:0] _io_rw_rdata_T_1 = decoded_1 ? _T_16 : 32'h0;
  wire [31:0] _io_rw_rdata_T_2 = decoded_2 ? reg_bp_0_address : 32'h0;
  wire [31:0] _io_rw_rdata_T_4 = decoded_4 ? reg_misa : 32'h0;
  wire [31:0] _io_rw_rdata_T_5 = decoded_5 ? read_mstatus : 32'h0;
  wire [31:0] _io_rw_rdata_T_6 = decoded_6 ? read_mtvec : 32'h0;
  wire [15:0] _io_rw_rdata_T_7 = decoded_7 ? read_mip : 16'h0;
  wire [31:0] _io_rw_rdata_T_8 = decoded_8 ? reg_mie : 32'h0;
  wire [31:0] _io_rw_rdata_T_9 = decoded_9 ? reg_mscratch : 32'h0;
  wire [31:0] _io_rw_rdata_T_10 = decoded_10 ? _T_22 : 32'h0;
  wire [31:0] _io_rw_rdata_T_11 = decoded_11 ? reg_mtval : 32'h0;
  wire [31:0] _io_rw_rdata_T_12 = decoded_12 ? reg_mcause : 32'h0;
  wire  _io_rw_rdata_T_13 = decoded_13 & io_hartid;
  wire [31:0] _io_rw_rdata_T_14 = decoded_14 ? _T_23 : 32'h0;
  wire [31:0] _io_rw_rdata_T_15 = decoded_15 ? _T_28 : 32'h0;
  wire [31:0] _io_rw_rdata_T_16 = decoded_16 ? reg_dscratch0 : 32'h0;
  wire [4:0] _io_rw_rdata_T_17 = decoded_17 ? reg_fflags : 5'h0;
  wire [2:0] _io_rw_rdata_T_18 = decoded_18 ? reg_frm : 3'h0;
  wire [7:0] _io_rw_rdata_T_19 = decoded_19 ? read_fcsr : 8'h0;
  wire [2:0] _io_rw_rdata_T_20 = decoded_20 ? reg_mcountinhibit : 3'h0;
  wire [63:0] _io_rw_rdata_T_21 = decoded_21 ? value_1 : 64'h0;
  wire [63:0] _io_rw_rdata_T_22 = decoded_22 ? value : 64'h0;
  wire [31:0] _io_rw_rdata_T_168 = decoded_168 ? read_mcounteren : 32'h0;
  wire [63:0] _io_rw_rdata_T_169 = decoded_169 ? value_1 : 64'h0;
  wire [63:0] _io_rw_rdata_T_170 = decoded_170 ? value : 64'h0;
  wire [31:0] _io_rw_rdata_T_171 = decoded_171 ? value_1[63:32] : 32'h0;
  wire [31:0] _io_rw_rdata_T_172 = decoded_172 ? value[63:32] : 32'h0;
  wire [31:0] _io_rw_rdata_T_173 = decoded_173 ? value_1[63:32] : 32'h0;
  wire [31:0] _io_rw_rdata_T_174 = decoded_174 ? value[63:32] : 32'h0;
  wire [31:0] _io_rw_rdata_T_175 = decoded_175 ? _T_91[31:0] : 32'h0;
  wire [31:0] _io_rw_rdata_T_176 = decoded_176 ? read_sip : 32'h0;
  wire [31:0] _io_rw_rdata_T_177 = decoded_177 ? read_sie : 32'h0;
  wire [31:0] _io_rw_rdata_T_178 = decoded_178 ? reg_sscratch : 32'h0;
  wire [31:0] _io_rw_rdata_T_179 = decoded_179 ? reg_scause : 32'h0;
  wire [31:0] _io_rw_rdata_T_180 = decoded_180 ? reg_stval : 32'h0;
  wire [31:0] _io_rw_rdata_T_181 = decoded_181 ? _T_93 : 32'h0;
  wire [31:0] _io_rw_rdata_T_182 = decoded_182 ? _T_98 : 32'h0;
  wire [31:0] _io_rw_rdata_T_183 = decoded_183 ? read_stvec : 32'h0;
  wire [31:0] _io_rw_rdata_T_184 = decoded_184 ? read_scounteren : 32'h0;
  wire [31:0] _io_rw_rdata_T_185 = decoded_185 ? read_mideleg : 32'h0;
  wire [31:0] _io_rw_rdata_T_186 = decoded_186 ? read_medeleg : 32'h0;
  wire [31:0] _io_rw_rdata_T_187 = decoded_187 ? _T_103 : 32'h0;
  wire [31:0] _io_rw_rdata_T_188 = decoded_188 ? _T_108 : 32'h0;
  wire [29:0] _io_rw_rdata_T_191 = decoded_191 ? reg_pmp_0_addr : 30'h0;
  wire [29:0] _io_rw_rdata_T_192 = decoded_192 ? reg_pmp_1_addr : 30'h0;
  wire [29:0] _io_rw_rdata_T_193 = decoded_193 ? reg_pmp_2_addr : 30'h0;
  wire [29:0] _io_rw_rdata_T_194 = decoded_194 ? reg_pmp_3_addr : 30'h0;
  wire [29:0] _io_rw_rdata_T_195 = decoded_195 ? reg_pmp_4_addr : 30'h0;
  wire [29:0] _io_rw_rdata_T_196 = decoded_196 ? reg_pmp_5_addr : 30'h0;
  wire [29:0] _io_rw_rdata_T_197 = decoded_197 ? reg_pmp_6_addr : 30'h0;
  wire [29:0] _io_rw_rdata_T_198 = decoded_198 ? reg_pmp_7_addr : 30'h0;
  wire [31:0] _io_rw_rdata_T_207 = decoded_207 ? reg_custom_0 : 32'h0;
  wire [31:0] _io_rw_rdata_T_208 = decoded_208 ? 32'h1 : 32'h0;
  wire [31:0] _io_rw_rdata_T_210 = decoded_210 ? 32'h20181004 : 32'h0;
  wire [31:0] _io_rw_rdata_T_212 = _io_rw_rdata_T_1 | _io_rw_rdata_T_2;
  wire [31:0] _io_rw_rdata_T_214 = _io_rw_rdata_T_212 | _io_rw_rdata_T_4;
  wire [31:0] _io_rw_rdata_T_215 = _io_rw_rdata_T_214 | _io_rw_rdata_T_5;
  wire [31:0] _io_rw_rdata_T_216 = _io_rw_rdata_T_215 | _io_rw_rdata_T_6;
  wire [31:0] _GEN_672 = {{16'd0}, _io_rw_rdata_T_7};
  wire [31:0] _io_rw_rdata_T_217 = _io_rw_rdata_T_216 | _GEN_672;
  wire [31:0] _io_rw_rdata_T_218 = _io_rw_rdata_T_217 | _io_rw_rdata_T_8;
  wire [31:0] _io_rw_rdata_T_219 = _io_rw_rdata_T_218 | _io_rw_rdata_T_9;
  wire [31:0] _io_rw_rdata_T_220 = _io_rw_rdata_T_219 | _io_rw_rdata_T_10;
  wire [31:0] _io_rw_rdata_T_221 = _io_rw_rdata_T_220 | _io_rw_rdata_T_11;
  wire [31:0] _io_rw_rdata_T_222 = _io_rw_rdata_T_221 | _io_rw_rdata_T_12;
  wire [31:0] _GEN_673 = {{31'd0}, _io_rw_rdata_T_13};
  wire [31:0] _io_rw_rdata_T_223 = _io_rw_rdata_T_222 | _GEN_673;
  wire [31:0] _io_rw_rdata_T_224 = _io_rw_rdata_T_223 | _io_rw_rdata_T_14;
  wire [31:0] _io_rw_rdata_T_225 = _io_rw_rdata_T_224 | _io_rw_rdata_T_15;
  wire [31:0] _io_rw_rdata_T_226 = _io_rw_rdata_T_225 | _io_rw_rdata_T_16;
  wire [31:0] _GEN_674 = {{27'd0}, _io_rw_rdata_T_17};
  wire [31:0] _io_rw_rdata_T_227 = _io_rw_rdata_T_226 | _GEN_674;
  wire [31:0] _GEN_675 = {{29'd0}, _io_rw_rdata_T_18};
  wire [31:0] _io_rw_rdata_T_228 = _io_rw_rdata_T_227 | _GEN_675;
  wire [31:0] _GEN_676 = {{24'd0}, _io_rw_rdata_T_19};
  wire [31:0] _io_rw_rdata_T_229 = _io_rw_rdata_T_228 | _GEN_676;
  wire [31:0] _GEN_677 = {{29'd0}, _io_rw_rdata_T_20};
  wire [31:0] _io_rw_rdata_T_230 = _io_rw_rdata_T_229 | _GEN_677;
  wire [63:0] _GEN_678 = {{32'd0}, _io_rw_rdata_T_230};
  wire [63:0] _io_rw_rdata_T_231 = _GEN_678 | _io_rw_rdata_T_21;
  wire [63:0] _io_rw_rdata_T_232 = _io_rw_rdata_T_231 | _io_rw_rdata_T_22;
  wire [63:0] _GEN_679 = {{32'd0}, _io_rw_rdata_T_168};
  wire [63:0] _io_rw_rdata_T_378 = _io_rw_rdata_T_232 | _GEN_679;
  wire [63:0] _io_rw_rdata_T_379 = _io_rw_rdata_T_378 | _io_rw_rdata_T_169;
  wire [63:0] _io_rw_rdata_T_380 = _io_rw_rdata_T_379 | _io_rw_rdata_T_170;
  wire [63:0] _GEN_680 = {{32'd0}, _io_rw_rdata_T_171};
  wire [63:0] _io_rw_rdata_T_381 = _io_rw_rdata_T_380 | _GEN_680;
  wire [63:0] _GEN_681 = {{32'd0}, _io_rw_rdata_T_172};
  wire [63:0] _io_rw_rdata_T_382 = _io_rw_rdata_T_381 | _GEN_681;
  wire [63:0] _GEN_682 = {{32'd0}, _io_rw_rdata_T_173};
  wire [63:0] _io_rw_rdata_T_383 = _io_rw_rdata_T_382 | _GEN_682;
  wire [63:0] _GEN_683 = {{32'd0}, _io_rw_rdata_T_174};
  wire [63:0] _io_rw_rdata_T_384 = _io_rw_rdata_T_383 | _GEN_683;
  wire [63:0] _GEN_684 = {{32'd0}, _io_rw_rdata_T_175};
  wire [63:0] _io_rw_rdata_T_385 = _io_rw_rdata_T_384 | _GEN_684;
  wire [63:0] _GEN_685 = {{32'd0}, _io_rw_rdata_T_176};
  wire [63:0] _io_rw_rdata_T_386 = _io_rw_rdata_T_385 | _GEN_685;
  wire [63:0] _GEN_686 = {{32'd0}, _io_rw_rdata_T_177};
  wire [63:0] _io_rw_rdata_T_387 = _io_rw_rdata_T_386 | _GEN_686;
  wire [63:0] _GEN_687 = {{32'd0}, _io_rw_rdata_T_178};
  wire [63:0] _io_rw_rdata_T_388 = _io_rw_rdata_T_387 | _GEN_687;
  wire [63:0] _GEN_688 = {{32'd0}, _io_rw_rdata_T_179};
  wire [63:0] _io_rw_rdata_T_389 = _io_rw_rdata_T_388 | _GEN_688;
  wire [63:0] _GEN_689 = {{32'd0}, _io_rw_rdata_T_180};
  wire [63:0] _io_rw_rdata_T_390 = _io_rw_rdata_T_389 | _GEN_689;
  wire [63:0] _GEN_690 = {{32'd0}, _io_rw_rdata_T_181};
  wire [63:0] _io_rw_rdata_T_391 = _io_rw_rdata_T_390 | _GEN_690;
  wire [63:0] _GEN_691 = {{32'd0}, _io_rw_rdata_T_182};
  wire [63:0] _io_rw_rdata_T_392 = _io_rw_rdata_T_391 | _GEN_691;
  wire [63:0] _GEN_692 = {{32'd0}, _io_rw_rdata_T_183};
  wire [63:0] _io_rw_rdata_T_393 = _io_rw_rdata_T_392 | _GEN_692;
  wire [63:0] _GEN_693 = {{32'd0}, _io_rw_rdata_T_184};
  wire [63:0] _io_rw_rdata_T_394 = _io_rw_rdata_T_393 | _GEN_693;
  wire [63:0] _GEN_694 = {{32'd0}, _io_rw_rdata_T_185};
  wire [63:0] _io_rw_rdata_T_395 = _io_rw_rdata_T_394 | _GEN_694;
  wire [63:0] _GEN_695 = {{32'd0}, _io_rw_rdata_T_186};
  wire [63:0] _io_rw_rdata_T_396 = _io_rw_rdata_T_395 | _GEN_695;
  wire [63:0] _GEN_696 = {{32'd0}, _io_rw_rdata_T_187};
  wire [63:0] _io_rw_rdata_T_397 = _io_rw_rdata_T_396 | _GEN_696;
  wire [63:0] _GEN_697 = {{32'd0}, _io_rw_rdata_T_188};
  wire [63:0] _io_rw_rdata_T_398 = _io_rw_rdata_T_397 | _GEN_697;
  wire [63:0] _GEN_698 = {{34'd0}, _io_rw_rdata_T_191};
  wire [63:0] _io_rw_rdata_T_401 = _io_rw_rdata_T_398 | _GEN_698;
  wire [63:0] _GEN_699 = {{34'd0}, _io_rw_rdata_T_192};
  wire [63:0] _io_rw_rdata_T_402 = _io_rw_rdata_T_401 | _GEN_699;
  wire [63:0] _GEN_700 = {{34'd0}, _io_rw_rdata_T_193};
  wire [63:0] _io_rw_rdata_T_403 = _io_rw_rdata_T_402 | _GEN_700;
  wire [63:0] _GEN_701 = {{34'd0}, _io_rw_rdata_T_194};
  wire [63:0] _io_rw_rdata_T_404 = _io_rw_rdata_T_403 | _GEN_701;
  wire [63:0] _GEN_702 = {{34'd0}, _io_rw_rdata_T_195};
  wire [63:0] _io_rw_rdata_T_405 = _io_rw_rdata_T_404 | _GEN_702;
  wire [63:0] _GEN_703 = {{34'd0}, _io_rw_rdata_T_196};
  wire [63:0] _io_rw_rdata_T_406 = _io_rw_rdata_T_405 | _GEN_703;
  wire [63:0] _GEN_704 = {{34'd0}, _io_rw_rdata_T_197};
  wire [63:0] _io_rw_rdata_T_407 = _io_rw_rdata_T_406 | _GEN_704;
  wire [63:0] _GEN_705 = {{34'd0}, _io_rw_rdata_T_198};
  wire [63:0] _io_rw_rdata_T_408 = _io_rw_rdata_T_407 | _GEN_705;
  wire [63:0] _GEN_706 = {{32'd0}, _io_rw_rdata_T_207};
  wire [63:0] _io_rw_rdata_T_417 = _io_rw_rdata_T_408 | _GEN_706;
  wire [63:0] _GEN_707 = {{32'd0}, _io_rw_rdata_T_208};
  wire [63:0] _io_rw_rdata_T_418 = _io_rw_rdata_T_417 | _GEN_707;
  wire [63:0] _GEN_708 = {{32'd0}, _io_rw_rdata_T_210};
  wire [63:0] _io_rw_rdata_T_420 = _io_rw_rdata_T_418 | _GEN_708;
  wire  _T_537 = io_rw_cmd == 3'h5;
  wire  _T_538 = io_rw_cmd == 3'h6;
  wire  _T_539 = io_rw_cmd == 3'h7;
  wire [4:0] _reg_fflags_T = reg_fflags | io_fcsr_flags_bits;
  wire [4:0] _GEN_282 = io_fcsr_flags_valid ? _reg_fflags_T : reg_fflags;
  wire  csr_wen = _T_538 | _T_539 | _T_537;
  wire [104:0] _new_mstatus_WIRE = {{73'd0}, wdata};
  wire  new_mstatus_sie = _new_mstatus_WIRE[1];
  wire  new_mstatus_mie = _new_mstatus_WIRE[3];
  wire  new_mstatus_spie = _new_mstatus_WIRE[5];
  wire  new_mstatus_mpie = _new_mstatus_WIRE[7];
  wire  new_mstatus_spp = _new_mstatus_WIRE[8];
  wire [1:0] new_mstatus_mpp = _new_mstatus_WIRE[12:11];
  wire [1:0] new_mstatus_fs = _new_mstatus_WIRE[14:13];
  wire  new_mstatus_mprv = _new_mstatus_WIRE[17];
  wire  new_mstatus_sum = _new_mstatus_WIRE[18];
  wire  new_mstatus_mxr = _new_mstatus_WIRE[19];
  wire  new_mstatus_tvm = _new_mstatus_WIRE[20];
  wire  new_mstatus_tw = _new_mstatus_WIRE[21];
  wire  new_mstatus_tsr = _new_mstatus_WIRE[22];
  wire  _reg_mstatus_fs_T = |new_mstatus_fs;
  wire [1:0] _reg_mstatus_fs_T_2 = _reg_mstatus_fs_T ? 2'h3 : 2'h0;
  wire [1:0] _GEN_288 = decoded_5 ? {{1'd0}, new_mstatus_spp} : _GEN_264;
  wire  f = wdata[5];
  wire [31:0] _reg_misa_T = ~wdata;
  wire  _reg_misa_T_1 = ~f;
  wire [3:0] _reg_misa_T_2 = {_reg_misa_T_1, 3'h0};
  wire [31:0] _GEN_709 = {{28'd0}, _reg_misa_T_2};
  wire [31:0] _reg_misa_T_3 = _reg_misa_T | _GEN_709;
  wire [31:0] _reg_misa_T_4 = ~_reg_misa_T_3;
  wire [31:0] _reg_misa_T_5 = _reg_misa_T_4 & 32'h1025;
  wire [31:0] _reg_misa_T_7 = reg_misa & 32'hffffefda;
  wire [31:0] _reg_misa_T_8 = _reg_misa_T_5 | _reg_misa_T_7;
  wire [15:0] _new_mip_T_2 = io_rw_cmd[1] ? _read_hvip_T : 16'h0;
  wire [31:0] _GEN_710 = {{16'd0}, _new_mip_T_2};
  wire [31:0] _new_mip_T_3 = _GEN_710 | io_rw_wdata;
  wire [31:0] _new_mip_T_8 = _new_mip_T_3 & _wdata_T_6;
  wire  new_mip_ssip = _new_mip_T_8[1];
  wire  new_mip_stip = _new_mip_T_8[5];
  wire  new_mip_seip = _new_mip_T_8[9];
  wire [31:0] _reg_mie_T = wdata & 32'haaa;
  wire [31:0] _reg_mepc_T_1 = _reg_misa_T | 32'h1;
  wire [31:0] _reg_mepc_T_2 = ~_reg_mepc_T_1;
  wire [31:0] _reg_mcause_T = wdata & 32'h8000000f;
  wire [31:0] _reg_mcountinhibit_T_1 = wdata & 32'hfffffffd;
  wire [31:0] _GEN_309 = decoded_20 ? _reg_mcountinhibit_T_1 : {{29'd0}, reg_mcountinhibit};
  wire [63:0] _T_2725 = {value_1[63:32],wdata};
  wire [63:0] _GEN_310 = decoded_21 ? _T_2725 : {{57'd0}, _GEN_2};
  wire [63:0] _T_2728 = {wdata,value_1[31:0]};
  wire [63:0] _GEN_312 = decoded_171 ? _T_2728 : _GEN_310;
  wire [63:0] _T_2730 = {value[63:32],wdata};
  wire [63:0] _GEN_314 = decoded_22 ? _T_2730 : {{57'd0}, _GEN_0};
  wire [63:0] _T_2733 = {wdata,value[31:0]};
  wire [63:0] _GEN_316 = decoded_172 ? _T_2733 : _GEN_314;
  wire [31:0] _GEN_319 = decoded_17 ? wdata : {{27'd0}, _GEN_282};
  wire [31:0] _GEN_321 = decoded_18 ? wdata : {{29'd0}, reg_frm};
  wire [31:0] _GEN_323 = decoded_19 ? wdata : _GEN_319;
  wire [31:0] _GEN_324 = decoded_19 ? {{5'd0}, wdata[31:5]} : _GEN_321;
  wire [1:0] new_dcsr_prv = wdata[1:0];
  wire  new_dcsr_ebreaku = wdata[12];
  wire  new_dcsr_ebreaks = wdata[13];
  wire  new_dcsr_ebreakm = wdata[15];
  wire [1:0] _GEN_334 = decoded_175 ? {{1'd0}, new_mstatus_spp} : _GEN_288;
  wire [31:0] _new_sip_T = ~read_mideleg;
  wire [31:0] _new_sip_T_1 = _GEN_41 & _new_sip_T;
  wire [31:0] _new_sip_T_2 = wdata & read_mideleg;
  wire [31:0] _new_sip_T_3 = _new_sip_T_1 | _new_sip_T_2;
  wire  new_sip_ssip = _new_sip_T_3[1];
  wire [21:0] new_satp_ppn = wdata[21:0];
  wire  new_satp_mode = wdata[31];
  wire  _T_2734 = ~new_satp_mode;
  wire  _T_2736 = _T_2734 | new_satp_mode;
  wire [31:0] _reg_mie_T_1 = ~sie_mask;
  wire [31:0] _reg_mie_T_2 = reg_mie & _reg_mie_T_1;
  wire [31:0] _reg_mie_T_3 = wdata & sie_mask;
  wire [31:0] _reg_mie_T_4 = _reg_mie_T_2 | _reg_mie_T_3;
  wire [31:0] _reg_scause_T = wdata & 32'h8000001f;
  wire [31:0] _newBPC_T_2 = io_rw_cmd[1] ? _T_16 : 32'h0;
  wire [31:0] _newBPC_T_3 = _newBPC_T_2 | io_rw_wdata;
  wire [31:0] _newBPC_T_8 = _newBPC_T_3 & _wdata_T_6;
  wire  newBPC_action = _newBPC_T_8[12];
  wire  newBPC_dmode = _newBPC_T_8[27];
  wire  dMode = newBPC_dmode & reg_debug;
  wire  _GEN_356 = dMode & newBPC_action;
  wire  newCfg_r = wdata[0];
  wire  newCfg_w = wdata[1];
  wire  newCfg_x = wdata[2];
  wire [1:0] newCfg_a = wdata[4:3];
  wire  newCfg_l = wdata[7];
  wire  _T_2754 = ~reg_pmp_1_cfg_a[1] & reg_pmp_1_cfg_a[0];
  wire  _T_2756 = reg_pmp_0_cfg_l | reg_pmp_1_cfg_l & _T_2754;
  wire [31:0] _GEN_427 = decoded_191 & ~_T_2756 ? wdata : {{2'd0}, reg_pmp_0_addr};
  wire  newCfg_1_r = wdata[8];
  wire  newCfg_1_w = wdata[9];
  wire  newCfg_1_x = wdata[10];
  wire [1:0] newCfg_1_a = wdata[12:11];
  wire  newCfg_1_l = wdata[15];
  wire  _T_2764 = ~reg_pmp_2_cfg_a[1] & reg_pmp_2_cfg_a[0];
  wire  _T_2766 = reg_pmp_1_cfg_l | reg_pmp_2_cfg_l & _T_2764;
  wire [31:0] _GEN_434 = decoded_192 & ~_T_2766 ? wdata : {{2'd0}, reg_pmp_1_addr};
  wire  newCfg_2_r = wdata[16];
  wire  newCfg_2_w = wdata[17];
  wire  newCfg_2_x = wdata[18];
  wire [1:0] newCfg_2_a = wdata[20:19];
  wire  newCfg_2_l = wdata[23];
  wire  _T_2774 = ~reg_pmp_3_cfg_a[1] & reg_pmp_3_cfg_a[0];
  wire  _T_2776 = reg_pmp_2_cfg_l | reg_pmp_3_cfg_l & _T_2774;
  wire [31:0] _GEN_441 = decoded_193 & ~_T_2776 ? wdata : {{2'd0}, reg_pmp_2_addr};
  wire  newCfg_3_r = wdata[24];
  wire  newCfg_3_w = wdata[25];
  wire  newCfg_3_x = wdata[26];
  wire [1:0] newCfg_3_a = wdata[28:27];
  wire  newCfg_3_l = wdata[31];
  wire  _T_2784 = ~reg_pmp_4_cfg_a[1] & reg_pmp_4_cfg_a[0];
  wire  _T_2786 = reg_pmp_3_cfg_l | reg_pmp_4_cfg_l & _T_2784;
  wire [31:0] _GEN_448 = decoded_194 & ~_T_2786 ? wdata : {{2'd0}, reg_pmp_3_addr};
  wire  _T_2794 = ~reg_pmp_5_cfg_a[1] & reg_pmp_5_cfg_a[0];
  wire  _T_2796 = reg_pmp_4_cfg_l | reg_pmp_5_cfg_l & _T_2794;
  wire [31:0] _GEN_455 = decoded_195 & ~_T_2796 ? wdata : {{2'd0}, reg_pmp_4_addr};
  wire  _T_2804 = ~reg_pmp_6_cfg_a[1] & reg_pmp_6_cfg_a[0];
  wire  _T_2806 = reg_pmp_5_cfg_l | reg_pmp_6_cfg_l & _T_2804;
  wire [31:0] _GEN_462 = decoded_196 & ~_T_2806 ? wdata : {{2'd0}, reg_pmp_5_addr};
  wire  _T_2814 = ~reg_pmp_7_cfg_a[1] & reg_pmp_7_cfg_a[0];
  wire  _T_2816 = reg_pmp_6_cfg_l | reg_pmp_7_cfg_l & _T_2814;
  wire [31:0] _GEN_469 = decoded_197 & ~_T_2816 ? wdata : {{2'd0}, reg_pmp_6_addr};
  wire  _T_2826 = reg_pmp_7_cfg_l | reg_pmp_7_cfg_l & _T_2814;
  wire [31:0] _GEN_476 = decoded_198 & ~_T_2826 ? wdata : {{2'd0}, reg_pmp_7_addr};
  wire [31:0] _reg_custom_0_T = wdata & 32'h208;
  wire [31:0] _reg_custom_0_T_2 = reg_custom_0 & 32'hfffffdf7;
  wire [31:0] _reg_custom_0_T_3 = _reg_custom_0_T | _reg_custom_0_T_2;
  wire [1:0] _GEN_489 = csr_wen ? _GEN_334 : _GEN_264;
  wire [31:0] _GEN_509 = csr_wen ? _GEN_309 : {{29'd0}, reg_mcountinhibit};
  wire [63:0] _GEN_510 = csr_wen ? _GEN_312 : {{57'd0}, _GEN_2};
  wire [63:0] _GEN_512 = csr_wen ? _GEN_316 : {{57'd0}, _GEN_0};
  wire [31:0] _GEN_515 = csr_wen ? _GEN_323 : {{27'd0}, _GEN_282};
  wire [31:0] _GEN_516 = csr_wen ? _GEN_324 : {{29'd0}, reg_frm};
  wire [31:0] _GEN_574 = csr_wen ? _GEN_427 : {{2'd0}, reg_pmp_0_addr};
  wire [31:0] _GEN_581 = csr_wen ? _GEN_434 : {{2'd0}, reg_pmp_1_addr};
  wire [31:0] _GEN_588 = csr_wen ? _GEN_441 : {{2'd0}, reg_pmp_2_addr};
  wire [31:0] _GEN_595 = csr_wen ? _GEN_448 : {{2'd0}, reg_pmp_3_addr};
  wire [31:0] _GEN_602 = csr_wen ? _GEN_455 : {{2'd0}, reg_pmp_4_addr};
  wire [31:0] _GEN_609 = csr_wen ? _GEN_462 : {{2'd0}, reg_pmp_5_addr};
  wire [31:0] _GEN_616 = csr_wen ? _GEN_469 : {{2'd0}, reg_pmp_6_addr};
  wire [31:0] _GEN_623 = csr_wen ? _GEN_476 : {{2'd0}, reg_pmp_7_addr};
  assign io_rw_rdata = _io_rw_rdata_T_420[31:0];
  assign io_decode_0_fp_illegal = io_status_fs == 2'h0 | ~reg_misa[5];
  assign io_decode_0_fp_csr = |_io_decode_0_fp_csr_T_1;
  assign io_decode_0_rocc_illegal = io_status_xs == 2'h0 | ~reg_misa[23];
  assign io_decode_0_read_illegal = _io_decode_0_read_illegal_T_17 | _io_decode_0_read_illegal_T_21;
  assign io_decode_0_write_illegal = &addr_1[11:10];
  assign io_decode_0_write_flush = ~(io_decode_0_write_flush_addr_m >= 12'h340 & io_decode_0_write_flush_addr_m <= 12'h343
    );
  assign io_decode_0_system_illegal = _io_decode_0_system_illegal_T_15 | _io_decode_0_system_illegal_T_18;
  assign io_csr_stall = reg_wfi | io_status_cease;
  assign io_eret = _exception_T | insn_ret;
  assign io_singleStep = reg_dcsr_step & _T_397;
  assign io_status_debug = reg_debug;
  assign io_status_cease = io_status_cease_r;
  assign io_status_wfi = reg_wfi;
  assign io_status_isa = reg_misa;
  assign io_status_dprv = reg_mstatus_mprv & _T_397 ? reg_mstatus_mpp : reg_mstatus_prv;
  assign io_status_dv = 1'h0;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_v = 1'h0;
  assign io_status_sd = &io_status_fs | &io_status_xs | &io_status_vs;
  assign io_status_zero2 = 23'h0;
  assign io_status_mpv = 1'h0;
  assign io_status_gva = reg_mstatus_gva;
  assign io_status_mbe = 1'h0;
  assign io_status_sbe = 1'h0;
  assign io_status_sxl = 2'h1;
  assign io_status_uxl = 2'h1;
  assign io_status_sd_rv32 = io_status_sd;
  assign io_status_zero1 = 8'h0;
  assign io_status_tsr = reg_mstatus_tsr;
  assign io_status_tw = reg_mstatus_tw;
  assign io_status_tvm = reg_mstatus_tvm;
  assign io_status_mxr = reg_mstatus_mxr;
  assign io_status_sum = reg_mstatus_sum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = 2'h0;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_vs = 2'h0;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_ube = 1'h0;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = 1'h0;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = 1'h0;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = 1'h0;
  assign io_ptbr_mode = reg_satp_mode;
  assign io_ptbr_ppn = reg_satp_ppn;
  assign io_evec = insn_ret ? _GEN_250 : tvec;
  assign io_time = value_1[31:0];
  assign io_fcsr_rm = reg_frm;
  assign io_interrupt = (anyInterrupt & ~io_singleStep | reg_singleStepped) & ~(reg_debug | io_status_cease);
  assign io_interrupt_cause = 32'h80000000 + _GEN_663;
  assign io_bp_0_control_action = reg_bp_0_control_action;
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch;
  assign io_bp_0_control_m = reg_bp_0_control_m;
  assign io_bp_0_control_s = reg_bp_0_control_s;
  assign io_bp_0_control_u = reg_bp_0_control_u;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_address = reg_bp_0_address;
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l;
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a;
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x;
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w;
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r;
  assign io_pmp_0_addr = reg_pmp_0_addr;
  assign io_pmp_0_mask = _pmp_mask_T_4[31:0];
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l;
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a;
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x;
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w;
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r;
  assign io_pmp_1_addr = reg_pmp_1_addr;
  assign io_pmp_1_mask = _pmp_mask_T_9[31:0];
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l;
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a;
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x;
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w;
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r;
  assign io_pmp_2_addr = reg_pmp_2_addr;
  assign io_pmp_2_mask = _pmp_mask_T_14[31:0];
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l;
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a;
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x;
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w;
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r;
  assign io_pmp_3_addr = reg_pmp_3_addr;
  assign io_pmp_3_mask = _pmp_mask_T_19[31:0];
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l;
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a;
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x;
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w;
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r;
  assign io_pmp_4_addr = reg_pmp_4_addr;
  assign io_pmp_4_mask = _pmp_mask_T_24[31:0];
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l;
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a;
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x;
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w;
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r;
  assign io_pmp_5_addr = reg_pmp_5_addr;
  assign io_pmp_5_mask = _pmp_mask_T_29[31:0];
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l;
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a;
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x;
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w;
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r;
  assign io_pmp_6_addr = reg_pmp_6_addr;
  assign io_pmp_6_mask = _pmp_mask_T_34[31:0];
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l;
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a;
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x;
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w;
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r;
  assign io_pmp_7_addr = reg_pmp_7_addr;
  assign io_pmp_7_mask = _pmp_mask_T_39[31:0];
  assign io_inhibit_cycle = reg_mcountinhibit[0];
  assign io_trace_0_valid = io_retire > 1'h0 | io_trace_0_exception;
  assign io_trace_0_iaddr = io_pc;
  assign io_trace_0_insn = io_inst_0;
  assign io_trace_0_exception = insn_call | insn_break | io_exception;
  assign io_customCSRs_0_value = reg_custom_0;
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if (new_prv == 2'h2) begin
      reg_mstatus_prv <= 2'h0;
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_mstatus_prv <= {{1'd0}, reg_mstatus_spp};
      end else begin
        reg_mstatus_prv <= _GEN_236;
      end
    end else if (exception) begin
      reg_mstatus_prv <= _GEN_150;
    end
    if (reset) begin
      reg_mstatus_gva <= 1'h0;
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (!(delegate)) begin
          reg_mstatus_gva <= io_gva;
        end
      end
    end
    if (reset) begin
      reg_mstatus_tsr <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_5) begin
        reg_mstatus_tsr <= new_mstatus_tsr;
      end
    end
    if (reset) begin
      reg_mstatus_tw <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_5) begin
        reg_mstatus_tw <= new_mstatus_tw;
      end
    end
    if (reset) begin
      reg_mstatus_tvm <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_5) begin
        reg_mstatus_tvm <= new_mstatus_tvm;
      end
    end
    if (reset) begin
      reg_mstatus_mxr <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_175) begin
        reg_mstatus_mxr <= new_mstatus_mxr;
      end else if (decoded_5) begin
        reg_mstatus_mxr <= new_mstatus_mxr;
      end
    end
    if (reset) begin
      reg_mstatus_sum <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_175) begin
        reg_mstatus_sum <= new_mstatus_sum;
      end else if (decoded_5) begin
        reg_mstatus_sum <= new_mstatus_sum;
      end
    end
    if (reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_5) begin
        reg_mstatus_mprv <= new_mstatus_mprv;
      end else begin
        reg_mstatus_mprv <= _GEN_278;
      end
    end else begin
      reg_mstatus_mprv <= _GEN_278;
    end
    if (reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_175) begin
        reg_mstatus_fs <= _reg_mstatus_fs_T_2;
      end else if (decoded_5) begin
        reg_mstatus_fs <= _reg_mstatus_fs_T_2;
      end
    end
    if (reset) begin
      reg_mstatus_mpp <= 2'h3;
    end else if (csr_wen) begin
      if (decoded_5) begin
        if (new_mstatus_mpp == 2'h2) begin
          reg_mstatus_mpp <= 2'h0;
        end else begin
          reg_mstatus_mpp <= new_mstatus_mpp;
        end
      end else begin
        reg_mstatus_mpp <= _GEN_275;
      end
    end else begin
      reg_mstatus_mpp <= _GEN_275;
    end
    if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_489[0];
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_5) begin
        reg_mstatus_mpie <= new_mstatus_mpie;
      end else begin
        reg_mstatus_mpie <= _GEN_274;
      end
    end else begin
      reg_mstatus_mpie <= _GEN_274;
    end
    if (reset) begin
      reg_mstatus_spie <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_175) begin
        reg_mstatus_spie <= new_mstatus_spie;
      end else if (decoded_5) begin
        reg_mstatus_spie <= new_mstatus_spie;
      end else begin
        reg_mstatus_spie <= _GEN_263;
      end
    end else begin
      reg_mstatus_spie <= _GEN_263;
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_5) begin
        reg_mstatus_mie <= new_mstatus_mie;
      end else begin
        reg_mstatus_mie <= _GEN_273;
      end
    end else begin
      reg_mstatus_mie <= _GEN_273;
    end
    if (reset) begin
      reg_mstatus_sie <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_175) begin
        reg_mstatus_sie <= new_mstatus_sie;
      end else if (decoded_5) begin
        reg_mstatus_sie <= new_mstatus_sie;
      end else begin
        reg_mstatus_sie <= _GEN_262;
      end
    end else begin
      reg_mstatus_sie <= _GEN_262;
    end
    if (reset) begin
      reg_dcsr_prv <= 2'h3;
    end else if (csr_wen) begin
      if (decoded_14) begin
        if (new_dcsr_prv == 2'h2) begin
          reg_dcsr_prv <= 2'h0;
        end else begin
          reg_dcsr_prv <= new_dcsr_prv;
        end
      end else begin
        reg_dcsr_prv <= _GEN_185;
      end
    end else begin
      reg_dcsr_prv <= _GEN_185;
    end
    if (_io_interrupt_T) begin
      reg_singleStepped <= 1'h0;
    end else begin
      reg_singleStepped <= _GEN_48;
    end
    if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_14) begin
        reg_dcsr_ebreakm <= new_dcsr_ebreakm;
      end
    end
    if (reset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_14) begin
        reg_dcsr_ebreaks <= new_dcsr_ebreaks;
      end
    end
    if (reset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_14) begin
        reg_dcsr_ebreaku <= new_dcsr_ebreaku;
      end
    end
    if (reset) begin
      reg_debug <= 1'h0;
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_debug <= _GEN_182;
      end else if (io_rw_addr[10] & io_rw_addr[7]) begin
        reg_debug <= 1'h0;
      end else begin
        reg_debug <= _GEN_182;
      end
    end else begin
      reg_debug <= _GEN_182;
    end
    if (csr_wen) begin
      if (decoded_185) begin
        reg_mideleg <= wdata;
      end
    end
    if (csr_wen) begin
      if (decoded_186) begin
        reg_medeleg <= wdata;
      end
    end
    if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          reg_dcsr_cause <= _reg_dcsr_cause_T_2;
        end
      end
    end
    if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_14) begin
        reg_dcsr_step <= wdata[2];
      end
    end
    if (csr_wen) begin
      if (decoded_15) begin
        reg_dpc <= _reg_mepc_T_2;
      end else begin
        reg_dpc <= _GEN_183;
      end
    end else begin
      reg_dpc <= _GEN_183;
    end
    if (csr_wen) begin
      if (decoded_16) begin
        reg_dscratch0 <= wdata;
      end
    end
    if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_dmode <= dMode;
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_action <= _GEN_356;
        end
      end
    end
    if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_tmatch <= wdata[8:7];
        end
      end
    end
    if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_m <= wdata[6];
        end
      end
    end
    if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_s <= wdata[4];
        end
      end
    end
    if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_u <= wdata[3];
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_x <= wdata[2];
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_w <= wdata[1];
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_1) begin
          reg_bp_0_control_r <= wdata[0];
        end
      end
    end
    if (csr_wen) begin
      if (~reg_bp_0_control_dmode | reg_debug) begin
        if (decoded_2) begin
          reg_bp_0_address <= wdata;
        end
      end
    end
    if (reset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_0_cfg_l) begin
        reg_pmp_0_cfg_l <= newCfg_l;
      end
    end
    if (reset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_0_cfg_l) begin
        reg_pmp_0_cfg_a <= newCfg_a;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_0_cfg_l) begin
        reg_pmp_0_cfg_x <= newCfg_x;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_0_cfg_l) begin
        reg_pmp_0_cfg_w <= newCfg_w & newCfg_r;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_0_cfg_l) begin
        reg_pmp_0_cfg_r <= newCfg_r;
      end
    end
    reg_pmp_0_addr <= _GEN_574[29:0];
    if (reset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_1_cfg_l) begin
        reg_pmp_1_cfg_l <= newCfg_1_l;
      end
    end
    if (reset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_1_cfg_l) begin
        reg_pmp_1_cfg_a <= newCfg_1_a;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_1_cfg_l) begin
        reg_pmp_1_cfg_x <= newCfg_1_x;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_1_cfg_l) begin
        reg_pmp_1_cfg_w <= newCfg_1_w & newCfg_1_r;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_1_cfg_l) begin
        reg_pmp_1_cfg_r <= newCfg_1_r;
      end
    end
    reg_pmp_1_addr <= _GEN_581[29:0];
    if (reset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_2_cfg_l) begin
        reg_pmp_2_cfg_l <= newCfg_2_l;
      end
    end
    if (reset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_2_cfg_l) begin
        reg_pmp_2_cfg_a <= newCfg_2_a;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_2_cfg_l) begin
        reg_pmp_2_cfg_x <= newCfg_2_x;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_2_cfg_l) begin
        reg_pmp_2_cfg_w <= newCfg_2_w & newCfg_2_r;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_2_cfg_l) begin
        reg_pmp_2_cfg_r <= newCfg_2_r;
      end
    end
    reg_pmp_2_addr <= _GEN_588[29:0];
    if (reset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_3_cfg_l) begin
        reg_pmp_3_cfg_l <= newCfg_3_l;
      end
    end
    if (reset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_3_cfg_l) begin
        reg_pmp_3_cfg_a <= newCfg_3_a;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_3_cfg_l) begin
        reg_pmp_3_cfg_x <= newCfg_3_x;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_3_cfg_l) begin
        reg_pmp_3_cfg_w <= newCfg_3_w & newCfg_3_r;
      end
    end
    if (csr_wen) begin
      if (decoded_187 & ~reg_pmp_3_cfg_l) begin
        reg_pmp_3_cfg_r <= newCfg_3_r;
      end
    end
    reg_pmp_3_addr <= _GEN_595[29:0];
    if (reset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_4_cfg_l) begin
        reg_pmp_4_cfg_l <= newCfg_l;
      end
    end
    if (reset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_4_cfg_l) begin
        reg_pmp_4_cfg_a <= newCfg_a;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_4_cfg_l) begin
        reg_pmp_4_cfg_x <= newCfg_x;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_4_cfg_l) begin
        reg_pmp_4_cfg_w <= newCfg_w & newCfg_r;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_4_cfg_l) begin
        reg_pmp_4_cfg_r <= newCfg_r;
      end
    end
    reg_pmp_4_addr <= _GEN_602[29:0];
    if (reset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_5_cfg_l) begin
        reg_pmp_5_cfg_l <= newCfg_1_l;
      end
    end
    if (reset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_5_cfg_l) begin
        reg_pmp_5_cfg_a <= newCfg_1_a;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_5_cfg_l) begin
        reg_pmp_5_cfg_x <= newCfg_1_x;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_5_cfg_l) begin
        reg_pmp_5_cfg_w <= newCfg_1_w & newCfg_1_r;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_5_cfg_l) begin
        reg_pmp_5_cfg_r <= newCfg_1_r;
      end
    end
    reg_pmp_5_addr <= _GEN_609[29:0];
    if (reset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_6_cfg_l) begin
        reg_pmp_6_cfg_l <= newCfg_2_l;
      end
    end
    if (reset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_6_cfg_l) begin
        reg_pmp_6_cfg_a <= newCfg_2_a;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_6_cfg_l) begin
        reg_pmp_6_cfg_x <= newCfg_2_x;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_6_cfg_l) begin
        reg_pmp_6_cfg_w <= newCfg_2_w & newCfg_2_r;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_6_cfg_l) begin
        reg_pmp_6_cfg_r <= newCfg_2_r;
      end
    end
    reg_pmp_6_addr <= _GEN_616[29:0];
    if (reset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_7_cfg_l) begin
        reg_pmp_7_cfg_l <= newCfg_3_l;
      end
    end
    if (reset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_7_cfg_l) begin
        reg_pmp_7_cfg_a <= newCfg_3_a;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_7_cfg_l) begin
        reg_pmp_7_cfg_x <= newCfg_3_x;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_7_cfg_l) begin
        reg_pmp_7_cfg_w <= newCfg_3_w & newCfg_3_r;
      end
    end
    if (csr_wen) begin
      if (decoded_188 & ~reg_pmp_7_cfg_l) begin
        reg_pmp_7_cfg_r <= newCfg_3_r;
      end
    end
    reg_pmp_7_addr <= _GEN_623[29:0];
    if (csr_wen) begin
      if (decoded_177) begin
        reg_mie <= _reg_mie_T_4;
      end else if (decoded_8) begin
        reg_mie <= _reg_mie_T;
      end
    end
    if (csr_wen) begin
      if (decoded_7) begin
        reg_mip_seip <= new_mip_seip;
      end
    end
    if (csr_wen) begin
      if (decoded_7) begin
        reg_mip_stip <= new_mip_stip;
      end
    end
    if (csr_wen) begin
      if (decoded_176) begin
        reg_mip_ssip <= new_sip_ssip;
      end else if (decoded_7) begin
        reg_mip_ssip <= new_mip_ssip;
      end
    end
    if (csr_wen) begin
      if (decoded_10) begin
        reg_mepc <= _reg_mepc_T_2;
      end else begin
        reg_mepc <= _GEN_211;
      end
    end else begin
      reg_mepc <= _GEN_211;
    end
    if (reset) begin
      reg_mcause <= 32'h0;
    end else if (csr_wen) begin
      if (decoded_12) begin
        reg_mcause <= _reg_mcause_T;
      end else begin
        reg_mcause <= _GEN_212;
      end
    end else begin
      reg_mcause <= _GEN_212;
    end
    if (csr_wen) begin
      if (decoded_11) begin
        reg_mtval <= wdata;
      end else begin
        reg_mtval <= _GEN_213;
      end
    end else begin
      reg_mtval <= _GEN_213;
    end
    if (csr_wen) begin
      if (decoded_9) begin
        reg_mscratch <= wdata;
      end
    end
    if (reset) begin
      reg_mtvec <= 32'h0;
    end else if (csr_wen) begin
      if (decoded_6) begin
        reg_mtvec <= wdata;
      end
    end
    if (csr_wen) begin
      if (decoded_168) begin
        reg_mcounteren <= wdata;
      end
    end
    if (csr_wen) begin
      if (decoded_184) begin
        reg_scounteren <= wdata;
      end
    end
    if (csr_wen) begin
      if (decoded_182) begin
        reg_sepc <= _reg_mepc_T_2;
      end else begin
        reg_sepc <= _GEN_202;
      end
    end else begin
      reg_sepc <= _GEN_202;
    end
    if (csr_wen) begin
      if (decoded_179) begin
        reg_scause <= _reg_scause_T;
      end else begin
        reg_scause <= _GEN_203;
      end
    end else begin
      reg_scause <= _GEN_203;
    end
    if (csr_wen) begin
      if (decoded_180) begin
        reg_stval <= wdata;
      end else begin
        reg_stval <= _GEN_204;
      end
    end else begin
      reg_stval <= _GEN_204;
    end
    if (csr_wen) begin
      if (decoded_178) begin
        reg_sscratch <= wdata;
      end
    end
    if (csr_wen) begin
      if (decoded_183) begin
        reg_stvec <= wdata;
      end
    end
    if (reset) begin
      reg_satp_mode <= 1'h0;
    end else if (csr_wen) begin
      if (decoded_181) begin
        if (_T_2736) begin
          reg_satp_mode <= new_satp_mode;
        end
      end
    end
    if (csr_wen) begin
      if (decoded_181) begin
        if (_T_2736) begin
          reg_satp_ppn <= {{2'd0}, new_satp_ppn[19:0]};
        end
      end
    end
    reg_fflags <= _GEN_515[4:0];
    reg_frm <= _GEN_516[2:0];
    if (reset) begin
      reg_mcountinhibit <= 3'h0;
    end else begin
      reg_mcountinhibit <= _GEN_509[2:0];
    end
    if (reset) begin
      small_ <= 6'h0;
    end else begin
      small_ <= _GEN_512[5:0];
    end
    if (reset) begin
      large_ <= 58'h0;
    end else if (csr_wen) begin
      if (decoded_172) begin
        large_ <= _T_2733[63:6];
      end else if (decoded_22) begin
        large_ <= _T_2730[63:6];
      end else begin
        large_ <= _GEN_1;
      end
    end else begin
      large_ <= _GEN_1;
    end
    if (reset) begin
      reg_misa <= 32'h40941125;
    end else if (csr_wen) begin
      if (decoded_4) begin
        if (~io_pc[1] | wdata[2]) begin
          reg_misa <= _reg_misa_T_8;
        end
      end
    end
    if (reset) begin
      reg_custom_0 <= 32'h208;
    end else if (csr_wen) begin
      if (decoded_207) begin
        reg_custom_0 <= _reg_custom_0_T_3;
      end
    end
    if (reset) begin
      io_status_cease_r <= 1'h0;
    end else begin
      io_status_cease_r <= _GEN_279;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_369 <= 3'h1) & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_369 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:957 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~reg_singleStepped | ~io_retire) & _T_373) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_373 & ~(~reg_singleStepped | ~io_retire)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CSR.scala:966 assert(!reg_singleStepped || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge io_ungated_clock) begin
    if (reset) begin
      reg_wfi <= 1'h0;
    end else if (|pending_interrupts | io_interrupts_debug | exception) begin
      reg_wfi <= 1'h0;
    end else begin
      reg_wfi <= _GEN_46;
    end
    if (reset) begin
      small_1 <= 6'h0;
    end else begin
      small_1 <= _GEN_510[5:0];
    end
    if (reset) begin
      large_1 <= 58'h0;
    end else if (csr_wen) begin
      if (decoded_171) begin
        large_1 <= _T_2728[63:6];
      end else if (decoded_21) begin
        large_1 <= _T_2725[63:6];
      end else begin
        large_1 <= _GEN_3;
      end
    end else begin
      large_1 <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_gva = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_tsr = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reg_mstatus_tw = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_mstatus_tvm = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_mstatus_mxr = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  reg_mstatus_sum = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  reg_mstatus_mprv = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reg_mstatus_fs = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reg_mstatus_mpp = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reg_mstatus_spp = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reg_mstatus_spie = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  reg_mstatus_sie = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_dcsr_prv = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  reg_singleStepped = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reg_dcsr_ebreaks = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  reg_dcsr_ebreaku = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  reg_debug = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  reg_mideleg = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_medeleg = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_dcsr_cause = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  reg_dpc = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_dscratch0 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_bp_0_control_dmode = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  reg_bp_0_control_action = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  reg_bp_0_control_tmatch = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  reg_bp_0_control_m = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  reg_bp_0_control_s = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  reg_bp_0_control_u = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  reg_bp_0_control_x = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  reg_bp_0_control_w = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  reg_bp_0_control_r = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  reg_bp_0_address = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  reg_pmp_0_cfg_l = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  reg_pmp_0_cfg_a = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  reg_pmp_0_cfg_x = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  reg_pmp_0_cfg_w = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  reg_pmp_0_cfg_r = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  reg_pmp_0_addr = _RAND_42[29:0];
  _RAND_43 = {1{`RANDOM}};
  reg_pmp_1_cfg_l = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  reg_pmp_1_cfg_a = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  reg_pmp_1_cfg_x = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  reg_pmp_1_cfg_w = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  reg_pmp_1_cfg_r = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  reg_pmp_1_addr = _RAND_48[29:0];
  _RAND_49 = {1{`RANDOM}};
  reg_pmp_2_cfg_l = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  reg_pmp_2_cfg_a = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  reg_pmp_2_cfg_x = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  reg_pmp_2_cfg_w = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  reg_pmp_2_cfg_r = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  reg_pmp_2_addr = _RAND_54[29:0];
  _RAND_55 = {1{`RANDOM}};
  reg_pmp_3_cfg_l = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  reg_pmp_3_cfg_a = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  reg_pmp_3_cfg_x = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  reg_pmp_3_cfg_w = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  reg_pmp_3_cfg_r = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  reg_pmp_3_addr = _RAND_60[29:0];
  _RAND_61 = {1{`RANDOM}};
  reg_pmp_4_cfg_l = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  reg_pmp_4_cfg_a = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  reg_pmp_4_cfg_x = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  reg_pmp_4_cfg_w = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  reg_pmp_4_cfg_r = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  reg_pmp_4_addr = _RAND_66[29:0];
  _RAND_67 = {1{`RANDOM}};
  reg_pmp_5_cfg_l = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  reg_pmp_5_cfg_a = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  reg_pmp_5_cfg_x = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  reg_pmp_5_cfg_w = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  reg_pmp_5_cfg_r = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  reg_pmp_5_addr = _RAND_72[29:0];
  _RAND_73 = {1{`RANDOM}};
  reg_pmp_6_cfg_l = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  reg_pmp_6_cfg_a = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  reg_pmp_6_cfg_x = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  reg_pmp_6_cfg_w = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  reg_pmp_6_cfg_r = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  reg_pmp_6_addr = _RAND_78[29:0];
  _RAND_79 = {1{`RANDOM}};
  reg_pmp_7_cfg_l = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  reg_pmp_7_cfg_a = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  reg_pmp_7_cfg_x = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  reg_pmp_7_cfg_w = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  reg_pmp_7_cfg_r = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  reg_pmp_7_addr = _RAND_84[29:0];
  _RAND_85 = {1{`RANDOM}};
  reg_mie = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  reg_mip_seip = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  reg_mip_stip = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  reg_mip_ssip = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  reg_mepc = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  reg_mcause = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  reg_mtval = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  reg_mscratch = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  reg_mtvec = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  reg_mcounteren = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  reg_scounteren = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  reg_sepc = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  reg_scause = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  reg_stval = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  reg_sscratch = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  reg_stvec = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  reg_satp_mode = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  reg_satp_ppn = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  reg_wfi = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  reg_fflags = _RAND_104[4:0];
  _RAND_105 = {1{`RANDOM}};
  reg_frm = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  reg_mcountinhibit = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  small_ = _RAND_107[5:0];
  _RAND_108 = {2{`RANDOM}};
  large_ = _RAND_108[57:0];
  _RAND_109 = {1{`RANDOM}};
  small_1 = _RAND_109[5:0];
  _RAND_110 = {2{`RANDOM}};
  large_1 = _RAND_110[57:0];
  _RAND_111 = {1{`RANDOM}};
  reg_misa = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  reg_custom_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  io_status_cease_r = _RAND_113[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule