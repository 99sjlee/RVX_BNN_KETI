// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************


`ifndef RVX_GDEF_001
`define RVX_GDEF_001

`define RVX_GDEF_324 3
`define RVX_GDEF_202 3

`define RVX_GDEF_022 0
`define RVX_GDEF_066 4

`define RVX_GDEF_179 1
`define RVX_GDEF_060 0
`define RVX_GDEF_280 1

`define RVX_GDEF_106(SOURCE,SIZE) (`RVX_GDEF_179+`RVX_GDEF_324+SOURCE+SIZE)

`endif
