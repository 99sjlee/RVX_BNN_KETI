// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef __ERVP_MMIOX1_MEMORYMAP_OFFSET_H__
`define __ERVP_MMIOX1_MEMORYMAP_OFFSET_H__

`define BW_MMAP_OFFSET_ERVP_MMIOX1 7
`define ERVP_MMIOX1_ADDR_INTERVAL 8
`define BW_UNUSED_ERVP_MMIOX1 3
`define NUM_ERVP_MMIOX1_SUBMODULE 1

`define MMAP_SUBOFFSET_MMIO_CORE_CONFIG_SAWD (32'h 0)
`define MMAP_SUBOFFSET_MMIO_CORE_STATUS_SAWD (32'h 8)
`define MMAP_SUBOFFSET_MMIO_CORE_CLEAR (32'h 10)
`define MMAP_SUBOFFSET_MMIO_LOG_FIFO_SAWD (32'h 18)
`define MMAP_SUBOFFSET_MMIO_INST_FIFO_SAWD (32'h 20)
`define MMAP_SUBOFFSET_MMIO_INST_STATUS (32'h 28)
`define MMAP_SUBOFFSET_MMIO_INPUT_FIFO_SAWD (32'h 30)
`define MMAP_SUBOFFSET_MMIO_OUTPUT_FIFO_SAWD (32'h 38)
`define MMAP_SUBOFFSET_MMIO_FIFO_STATUS (32'h 40)
`define MMAP_SUBOFFSET_MMIO_ITR_REQUEST (32'h 48)
`define MMAP_SUBOFFSET_MMIO_ITR_STATUS (32'h 50)

`define MMAP_OFFSET_MMIO_CORE_CONFIG_SAWD (`MMAP_SUBOFFSET_MMIO_CORE_CONFIG_SAWD)
`define MMAP_OFFSET_MMIO_CORE_STATUS_SAWD (`MMAP_SUBOFFSET_MMIO_CORE_STATUS_SAWD)
`define MMAP_OFFSET_MMIO_CORE_CLEAR (`MMAP_SUBOFFSET_MMIO_CORE_CLEAR)
`define MMAP_OFFSET_MMIO_LOG_FIFO_SAWD (`MMAP_SUBOFFSET_MMIO_LOG_FIFO_SAWD)
`define MMAP_OFFSET_MMIO_INST_FIFO_SAWD (`MMAP_SUBOFFSET_MMIO_INST_FIFO_SAWD)
`define MMAP_OFFSET_MMIO_INST_STATUS (`MMAP_SUBOFFSET_MMIO_INST_STATUS)
`define MMAP_OFFSET_MMIO_INPUT_FIFO_SAWD (`MMAP_SUBOFFSET_MMIO_INPUT_FIFO_SAWD)
`define MMAP_OFFSET_MMIO_OUTPUT_FIFO_SAWD (`MMAP_SUBOFFSET_MMIO_OUTPUT_FIFO_SAWD)
`define MMAP_OFFSET_MMIO_FIFO_STATUS (`MMAP_SUBOFFSET_MMIO_FIFO_STATUS)
`define MMAP_OFFSET_MMIO_ITR_REQUEST (`MMAP_SUBOFFSET_MMIO_ITR_REQUEST)
`define MMAP_OFFSET_MMIO_ITR_STATUS (`MMAP_SUBOFFSET_MMIO_ITR_STATUS)

`define BW_MMIO_INST_STATUS 32
`define MMIO_INST_STATUS_DEFAULT_VALUE 0
`define MMIO_INST_STATUS_NUM_INFO_000 1
`define MMIO_INST_STATUS_NUM_INFO_001 2
`define MMIO_INST_STATUS_NUM_INFO_002 4
`define MMIO_INST_STATUS_NUM_INFO_003 8
`define MMIO_INST_STATUS_NUM_INFO_004 16
`define MMIO_INST_STATUS_NUM_INFO_005 32
`define MMIO_INST_STATUS_NUM_INFO_006 64
`define MMIO_INST_STATUS_NUM_INFO_007 128
`define MMIO_INST_STATUS_NUM_BUSY_000 256
`define MMIO_INST_STATUS_NUM_BUSY_001 512
`define MMIO_INST_STATUS_NUM_BUSY_002 1024
`define MMIO_INST_STATUS_NUM_BUSY_003 2048
`define MMIO_INST_STATUS_NUM_BUSY_004 4096
`define MMIO_INST_STATUS_NUM_BUSY_005 8192
`define MMIO_INST_STATUS_NUM_BUSY_006 16384
`define MMIO_INST_STATUS_NUM_BUSY_007 32768
`define MMIO_INST_STATUS_HAS_LOG 65536
`define MMIO_INST_STATUS_INDEX_NUM_INFO_000 0
`define MMIO_INST_STATUS_INDEX_NUM_INFO_001 1
`define MMIO_INST_STATUS_INDEX_NUM_INFO_002 2
`define MMIO_INST_STATUS_INDEX_NUM_INFO_003 3
`define MMIO_INST_STATUS_INDEX_NUM_INFO_004 4
`define MMIO_INST_STATUS_INDEX_NUM_INFO_005 5
`define MMIO_INST_STATUS_INDEX_NUM_INFO_006 6
`define MMIO_INST_STATUS_INDEX_NUM_INFO_007 7
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_000 8
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_001 9
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_002 10
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_003 11
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_004 12
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_005 13
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_006 14
`define MMIO_INST_STATUS_INDEX_NUM_BUSY_007 15
`define MMIO_INST_STATUS_INDEX_HAS_LOG 16
`define MMIO_INST_STATUS_NONE 0

`define BW_MMIO_CORE_CONFIG_SAWD 32
`define MMIO_CORE_CONFIG_SAWD_DEFAULT_VALUE 0

`define BW_MMIO_CORE_STATUS_SAWD 32
`define MMIO_CORE_STATUS_SAWD_DEFAULT_VALUE 0

`define BW_MMIO_CORE_CLEAR 1
`define MMIO_CORE_CLEAR_DEFAULT_VALUE 0

`define BW_MMIO_LOG_FIFO_SAWD 32
`define MMIO_LOG_FIFO_SAWD_DEFAULT_VALUE 0

`define BW_MMIO_INST_FIFO_SAWD 32
`define MMIO_INST_FIFO_SAWD_DEFAULT_VALUE 0

`define BW_MMIO_INPUT_FIFO_SAWD 32
`define MMIO_INPUT_FIFO_SAWD_DEFAULT_VALUE 0

`define BW_MMIO_OUTPUT_FIFO_SAWD 32
`define MMIO_OUTPUT_FIFO_SAWD_DEFAULT_VALUE 0

`define BW_MMIO_FIFO_STATUS 32
`define MMIO_FIFO_STATUS_DEFAULT_VALUE 0

`define BW_MMIO_ITR_REQUEST 32
`define MMIO_ITR_REQUEST_DEFAULT_VALUE 0

`define BW_MMIO_ITR_STATUS 32
`define MMIO_ITR_STATUS_DEFAULT_VALUE 0

`endif