// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_305
`define RVX_GDEF_305

`define RVX_GDEF_175 15
`define RVX_GDEF_112 8
`define RVX_GDEF_067 3
`define RVX_GDEF_216 5
`define RVX_GDEF_154 3
`define RVX_GDEF_071 0
`define RVX_GDEF_057 (32'h 0)
`define RVX_GDEF_096 1
`define RVX_GDEF_190 (32'h 1000)
`define RVX_GDEF_267 2
`define RVX_GDEF_069 (32'h 2000)
`define RVX_GDEF_276 3
`define RVX_GDEF_325 (32'h 3000)
`define RVX_GDEF_306 4
`define RVX_GDEF_346 (32'h 4000)

`define RVX_GDEF_213 8
`define RVX_GDEF_102 3

`define RVX_GDEF_055 5
`define RVX_GDEF_238 3
`define RVX_GDEF_416 (32'h 0)
`define RVX_GDEF_131 (32'h 8)
`define RVX_GDEF_050 (32'h 10)

`define RVX_GDEF_334 (`RVX_GDEF_190+`RVX_GDEF_416)
`define RVX_GDEF_013 (`RVX_GDEF_190+`RVX_GDEF_131)
`define RVX_GDEF_418 (`RVX_GDEF_190+`RVX_GDEF_050)

`define RVX_GDEF_161 12
`define RVX_GDEF_359 3

`define RVX_GDEF_429 10
`define RVX_GDEF_074 3

`define RVX_GDEF_200 10
`define RVX_GDEF_114 3

`define RVX_GDEF_412 8
`define RVX_GDEF_333 0

`define RVX_GDEF_002 8
`define RVX_GDEF_160 0

`define RVX_GDEF_100 1
`define RVX_GDEF_420 0

`endif