`default_nettype wire
module DCache(
  input         clock,
  input         reset,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output        auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [3:0]  auto_out_a_bits_mask,
  output [31:0] auto_out_a_bits_data,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output [31:0] auto_out_c_bits_address,
  output [31:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input         auto_out_d_bits_source,
  input  [2:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [31:0] auto_out_d_bits_data,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [2:0]  auto_out_e_bits_sink,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [6:0]  io_cpu_req_bits_tag,
  input  [4:0]  io_cpu_req_bits_cmd,
  input  [1:0]  io_cpu_req_bits_size,
  input         io_cpu_req_bits_signed,
  input  [1:0]  io_cpu_req_bits_dprv,
  input         io_cpu_req_bits_phys,
  input         io_cpu_s1_kill,
  input  [31:0] io_cpu_s1_data_data,
  input  [3:0]  io_cpu_s1_data_mask,
  output        io_cpu_s2_nack,
  output        io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_addr,
  output [6:0]  io_cpu_resp_bits_tag,
  output [4:0]  io_cpu_resp_bits_cmd,
  output [1:0]  io_cpu_resp_bits_size,
  output        io_cpu_resp_bits_signed,
  output [1:0]  io_cpu_resp_bits_dprv,
  output        io_cpu_resp_bits_dv,
  output [31:0] io_cpu_resp_bits_data,
  output [3:0]  io_cpu_resp_bits_mask,
  output        io_cpu_resp_bits_replay,
  output        io_cpu_resp_bits_has_data,
  output [31:0] io_cpu_resp_bits_data_word_bypass,
  output [31:0] io_cpu_resp_bits_data_raw,
  output [31:0] io_cpu_resp_bits_store_data,
  output        io_cpu_replay_next,
  output        io_cpu_s2_xcpt_ma_ld,
  output        io_cpu_s2_xcpt_ma_st,
  output        io_cpu_s2_xcpt_pf_ld,
  output        io_cpu_s2_xcpt_pf_st,
  output        io_cpu_s2_xcpt_gf_ld,
  output        io_cpu_s2_xcpt_gf_st,
  output        io_cpu_s2_xcpt_ae_ld,
  output        io_cpu_s2_xcpt_ae_st,
  output        io_cpu_ordered,
  output        io_cpu_perf_release,
  output        io_cpu_perf_grant,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [19:0] io_ptw_req_bits_bits_addr,
  output        io_ptw_req_bits_bits_need_gpa,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae_ptw,
  input         io_ptw_resp_bits_ae_final,
  input         io_ptw_resp_bits_pf,
  input  [43:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input         io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input         io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [31:0] tlb_io_req_bits_vaddr;
  wire  tlb_io_req_bits_passthrough;
  wire [1:0] tlb_io_req_bits_size;
  wire [4:0] tlb_io_req_bits_cmd;
  wire [1:0] tlb_io_req_bits_prv;
  wire  tlb_io_resp_miss;
  wire [31:0] tlb_io_resp_paddr;
  wire  tlb_io_resp_pf_ld;
  wire  tlb_io_resp_pf_st;
  wire  tlb_io_resp_ae_ld;
  wire  tlb_io_resp_ae_st;
  wire  tlb_io_resp_ma_ld;
  wire  tlb_io_resp_ma_st;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_sfence_valid;
  wire  tlb_io_sfence_bits_rs1;
  wire  tlb_io_sfence_bits_rs2;
  wire [31:0] tlb_io_sfence_bits_addr;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [19:0] tlb_io_ptw_req_bits_bits_addr;
  wire  tlb_io_ptw_req_bits_bits_need_gpa;
  wire  tlb_io_ptw_resp_valid;
  wire  tlb_io_ptw_resp_bits_ae_ptw;
  wire  tlb_io_ptw_resp_bits_ae_final;
  wire  tlb_io_ptw_resp_bits_pf;
  wire [43:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_a;
  wire  tlb_io_ptw_resp_bits_pte_g;
  wire  tlb_io_ptw_resp_bits_pte_u;
  wire  tlb_io_ptw_resp_bits_pte_x;
  wire  tlb_io_ptw_resp_bits_pte_w;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire  tlb_io_ptw_resp_bits_level;
  wire  tlb_io_ptw_resp_bits_homogeneous;
  wire  tlb_io_ptw_ptbr_mode;
  wire  tlb_io_ptw_status_debug;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_sum;
  wire  tlb_io_ptw_pmp_0_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a;
  wire  tlb_io_ptw_pmp_0_cfg_x;
  wire  tlb_io_ptw_pmp_0_cfg_w;
  wire  tlb_io_ptw_pmp_0_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_0_addr;
  wire [31:0] tlb_io_ptw_pmp_0_mask;
  wire  tlb_io_ptw_pmp_1_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a;
  wire  tlb_io_ptw_pmp_1_cfg_x;
  wire  tlb_io_ptw_pmp_1_cfg_w;
  wire  tlb_io_ptw_pmp_1_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_1_addr;
  wire [31:0] tlb_io_ptw_pmp_1_mask;
  wire  tlb_io_ptw_pmp_2_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a;
  wire  tlb_io_ptw_pmp_2_cfg_x;
  wire  tlb_io_ptw_pmp_2_cfg_w;
  wire  tlb_io_ptw_pmp_2_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_2_addr;
  wire [31:0] tlb_io_ptw_pmp_2_mask;
  wire  tlb_io_ptw_pmp_3_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a;
  wire  tlb_io_ptw_pmp_3_cfg_x;
  wire  tlb_io_ptw_pmp_3_cfg_w;
  wire  tlb_io_ptw_pmp_3_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_3_addr;
  wire [31:0] tlb_io_ptw_pmp_3_mask;
  wire  tlb_io_ptw_pmp_4_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a;
  wire  tlb_io_ptw_pmp_4_cfg_x;
  wire  tlb_io_ptw_pmp_4_cfg_w;
  wire  tlb_io_ptw_pmp_4_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_4_addr;
  wire [31:0] tlb_io_ptw_pmp_4_mask;
  wire  tlb_io_ptw_pmp_5_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a;
  wire  tlb_io_ptw_pmp_5_cfg_x;
  wire  tlb_io_ptw_pmp_5_cfg_w;
  wire  tlb_io_ptw_pmp_5_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_5_addr;
  wire [31:0] tlb_io_ptw_pmp_5_mask;
  wire  tlb_io_ptw_pmp_6_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a;
  wire  tlb_io_ptw_pmp_6_cfg_x;
  wire  tlb_io_ptw_pmp_6_cfg_w;
  wire  tlb_io_ptw_pmp_6_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_6_addr;
  wire [31:0] tlb_io_ptw_pmp_6_mask;
  wire  tlb_io_ptw_pmp_7_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a;
  wire  tlb_io_ptw_pmp_7_cfg_x;
  wire  tlb_io_ptw_pmp_7_cfg_w;
  wire  tlb_io_ptw_pmp_7_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_7_addr;
  wire [31:0] tlb_io_ptw_pmp_7_mask;
  wire [19:0] tlb_mpu_ppn_barrier_io_x_ppn;
  wire  tlb_mpu_ppn_barrier_io_x_u;
  wire  tlb_mpu_ppn_barrier_io_x_ae_ptw;
  wire  tlb_mpu_ppn_barrier_io_x_ae_final;
  wire  tlb_mpu_ppn_barrier_io_x_pf;
  wire  tlb_mpu_ppn_barrier_io_x_gf;
  wire  tlb_mpu_ppn_barrier_io_x_sw;
  wire  tlb_mpu_ppn_barrier_io_x_sx;
  wire  tlb_mpu_ppn_barrier_io_x_sr;
  wire  tlb_mpu_ppn_barrier_io_x_pw;
  wire  tlb_mpu_ppn_barrier_io_x_px;
  wire  tlb_mpu_ppn_barrier_io_x_pr;
  wire  tlb_mpu_ppn_barrier_io_x_ppp;
  wire  tlb_mpu_ppn_barrier_io_x_pal;
  wire  tlb_mpu_ppn_barrier_io_x_paa;
  wire  tlb_mpu_ppn_barrier_io_x_eff;
  wire  tlb_mpu_ppn_barrier_io_x_c;
  wire [19:0] tlb_mpu_ppn_barrier_io_y_ppn;
  wire  tlb_mpu_ppn_barrier_io_y_u;
  wire  tlb_mpu_ppn_barrier_io_y_ae_ptw;
  wire  tlb_mpu_ppn_barrier_io_y_ae_final;
  wire  tlb_mpu_ppn_barrier_io_y_pf;
  wire  tlb_mpu_ppn_barrier_io_y_gf;
  wire  tlb_mpu_ppn_barrier_io_y_sw;
  wire  tlb_mpu_ppn_barrier_io_y_sx;
  wire  tlb_mpu_ppn_barrier_io_y_sr;
  wire  tlb_mpu_ppn_barrier_io_y_pw;
  wire  tlb_mpu_ppn_barrier_io_y_px;
  wire  tlb_mpu_ppn_barrier_io_y_pr;
  wire  tlb_mpu_ppn_barrier_io_y_ppp;
  wire  tlb_mpu_ppn_barrier_io_y_pal;
  wire  tlb_mpu_ppn_barrier_io_y_paa;
  wire  tlb_mpu_ppn_barrier_io_y_eff;
  wire  tlb_mpu_ppn_barrier_io_y_c;
  wire [1:0] tlb_pmp_io_prv;
  wire  tlb_pmp_io_pmp_0_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_0_cfg_a;
  wire  tlb_pmp_io_pmp_0_cfg_x;
  wire  tlb_pmp_io_pmp_0_cfg_w;
  wire  tlb_pmp_io_pmp_0_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_0_addr;
  wire [31:0] tlb_pmp_io_pmp_0_mask;
  wire  tlb_pmp_io_pmp_1_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_1_cfg_a;
  wire  tlb_pmp_io_pmp_1_cfg_x;
  wire  tlb_pmp_io_pmp_1_cfg_w;
  wire  tlb_pmp_io_pmp_1_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_1_addr;
  wire [31:0] tlb_pmp_io_pmp_1_mask;
  wire  tlb_pmp_io_pmp_2_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_2_cfg_a;
  wire  tlb_pmp_io_pmp_2_cfg_x;
  wire  tlb_pmp_io_pmp_2_cfg_w;
  wire  tlb_pmp_io_pmp_2_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_2_addr;
  wire [31:0] tlb_pmp_io_pmp_2_mask;
  wire  tlb_pmp_io_pmp_3_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_3_cfg_a;
  wire  tlb_pmp_io_pmp_3_cfg_x;
  wire  tlb_pmp_io_pmp_3_cfg_w;
  wire  tlb_pmp_io_pmp_3_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_3_addr;
  wire [31:0] tlb_pmp_io_pmp_3_mask;
  wire  tlb_pmp_io_pmp_4_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_4_cfg_a;
  wire  tlb_pmp_io_pmp_4_cfg_x;
  wire  tlb_pmp_io_pmp_4_cfg_w;
  wire  tlb_pmp_io_pmp_4_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_4_addr;
  wire [31:0] tlb_pmp_io_pmp_4_mask;
  wire  tlb_pmp_io_pmp_5_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_5_cfg_a;
  wire  tlb_pmp_io_pmp_5_cfg_x;
  wire  tlb_pmp_io_pmp_5_cfg_w;
  wire  tlb_pmp_io_pmp_5_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_5_addr;
  wire [31:0] tlb_pmp_io_pmp_5_mask;
  wire  tlb_pmp_io_pmp_6_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_6_cfg_a;
  wire  tlb_pmp_io_pmp_6_cfg_x;
  wire  tlb_pmp_io_pmp_6_cfg_w;
  wire  tlb_pmp_io_pmp_6_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_6_addr;
  wire [31:0] tlb_pmp_io_pmp_6_mask;
  wire  tlb_pmp_io_pmp_7_cfg_l;
  wire [1:0] tlb_pmp_io_pmp_7_cfg_a;
  wire  tlb_pmp_io_pmp_7_cfg_x;
  wire  tlb_pmp_io_pmp_7_cfg_w;
  wire  tlb_pmp_io_pmp_7_cfg_r;
  wire [29:0] tlb_pmp_io_pmp_7_addr;
  wire [31:0] tlb_pmp_io_pmp_7_mask;
  wire [31:0] tlb_pmp_io_addr;
  wire  tlb_pmp_io_r;
  wire  tlb_pmp_io_w;
  wire  tlb_pmp_io_x;
  wire [19:0] tlb_entries_barrier_io_x_ppn;
  wire  tlb_entries_barrier_io_x_u;
  wire  tlb_entries_barrier_io_x_ae_ptw;
  wire  tlb_entries_barrier_io_x_ae_final;
  wire  tlb_entries_barrier_io_x_pf;
  wire  tlb_entries_barrier_io_x_gf;
  wire  tlb_entries_barrier_io_x_sw;
  wire  tlb_entries_barrier_io_x_sx;
  wire  tlb_entries_barrier_io_x_sr;
  wire  tlb_entries_barrier_io_x_pw;
  wire  tlb_entries_barrier_io_x_px;
  wire  tlb_entries_barrier_io_x_pr;
  wire  tlb_entries_barrier_io_x_ppp;
  wire  tlb_entries_barrier_io_x_pal;
  wire  tlb_entries_barrier_io_x_paa;
  wire  tlb_entries_barrier_io_x_eff;
  wire  tlb_entries_barrier_io_x_c;
  wire [19:0] tlb_entries_barrier_io_y_ppn;
  wire  tlb_entries_barrier_io_y_u;
  wire  tlb_entries_barrier_io_y_ae_ptw;
  wire  tlb_entries_barrier_io_y_ae_final;
  wire  tlb_entries_barrier_io_y_pf;
  wire  tlb_entries_barrier_io_y_gf;
  wire  tlb_entries_barrier_io_y_sw;
  wire  tlb_entries_barrier_io_y_sx;
  wire  tlb_entries_barrier_io_y_sr;
  wire  tlb_entries_barrier_io_y_pw;
  wire  tlb_entries_barrier_io_y_px;
  wire  tlb_entries_barrier_io_y_pr;
  wire  tlb_entries_barrier_io_y_ppp;
  wire  tlb_entries_barrier_io_y_pal;
  wire  tlb_entries_barrier_io_y_paa;
  wire  tlb_entries_barrier_io_y_eff;
  wire  tlb_entries_barrier_io_y_c;
  wire [19:0] tlb_entries_barrier_1_io_x_ppn;
  wire  tlb_entries_barrier_1_io_x_u;
  wire  tlb_entries_barrier_1_io_x_ae_ptw;
  wire  tlb_entries_barrier_1_io_x_ae_final;
  wire  tlb_entries_barrier_1_io_x_pf;
  wire  tlb_entries_barrier_1_io_x_gf;
  wire  tlb_entries_barrier_1_io_x_sw;
  wire  tlb_entries_barrier_1_io_x_sx;
  wire  tlb_entries_barrier_1_io_x_sr;
  wire  tlb_entries_barrier_1_io_x_pw;
  wire  tlb_entries_barrier_1_io_x_px;
  wire  tlb_entries_barrier_1_io_x_pr;
  wire  tlb_entries_barrier_1_io_x_ppp;
  wire  tlb_entries_barrier_1_io_x_pal;
  wire  tlb_entries_barrier_1_io_x_paa;
  wire  tlb_entries_barrier_1_io_x_eff;
  wire  tlb_entries_barrier_1_io_x_c;
  wire [19:0] tlb_entries_barrier_1_io_y_ppn;
  wire  tlb_entries_barrier_1_io_y_u;
  wire  tlb_entries_barrier_1_io_y_ae_ptw;
  wire  tlb_entries_barrier_1_io_y_ae_final;
  wire  tlb_entries_barrier_1_io_y_pf;
  wire  tlb_entries_barrier_1_io_y_gf;
  wire  tlb_entries_barrier_1_io_y_sw;
  wire  tlb_entries_barrier_1_io_y_sx;
  wire  tlb_entries_barrier_1_io_y_sr;
  wire  tlb_entries_barrier_1_io_y_pw;
  wire  tlb_entries_barrier_1_io_y_px;
  wire  tlb_entries_barrier_1_io_y_pr;
  wire  tlb_entries_barrier_1_io_y_ppp;
  wire  tlb_entries_barrier_1_io_y_pal;
  wire  tlb_entries_barrier_1_io_y_paa;
  wire  tlb_entries_barrier_1_io_y_eff;
  wire  tlb_entries_barrier_1_io_y_c;
  wire [19:0] tlb_entries_barrier_2_io_x_ppn;
  wire  tlb_entries_barrier_2_io_x_u;
  wire  tlb_entries_barrier_2_io_x_ae_ptw;
  wire  tlb_entries_barrier_2_io_x_ae_final;
  wire  tlb_entries_barrier_2_io_x_pf;
  wire  tlb_entries_barrier_2_io_x_gf;
  wire  tlb_entries_barrier_2_io_x_sw;
  wire  tlb_entries_barrier_2_io_x_sx;
  wire  tlb_entries_barrier_2_io_x_sr;
  wire  tlb_entries_barrier_2_io_x_pw;
  wire  tlb_entries_barrier_2_io_x_px;
  wire  tlb_entries_barrier_2_io_x_pr;
  wire  tlb_entries_barrier_2_io_x_ppp;
  wire  tlb_entries_barrier_2_io_x_pal;
  wire  tlb_entries_barrier_2_io_x_paa;
  wire  tlb_entries_barrier_2_io_x_eff;
  wire  tlb_entries_barrier_2_io_x_c;
  wire [19:0] tlb_entries_barrier_2_io_y_ppn;
  wire  tlb_entries_barrier_2_io_y_u;
  wire  tlb_entries_barrier_2_io_y_ae_ptw;
  wire  tlb_entries_barrier_2_io_y_ae_final;
  wire  tlb_entries_barrier_2_io_y_pf;
  wire  tlb_entries_barrier_2_io_y_gf;
  wire  tlb_entries_barrier_2_io_y_sw;
  wire  tlb_entries_barrier_2_io_y_sx;
  wire  tlb_entries_barrier_2_io_y_sr;
  wire  tlb_entries_barrier_2_io_y_pw;
  wire  tlb_entries_barrier_2_io_y_px;
  wire  tlb_entries_barrier_2_io_y_pr;
  wire  tlb_entries_barrier_2_io_y_ppp;
  wire  tlb_entries_barrier_2_io_y_pal;
  wire  tlb_entries_barrier_2_io_y_paa;
  wire  tlb_entries_barrier_2_io_y_eff;
  wire  tlb_entries_barrier_2_io_y_c;
  wire [19:0] tlb_entries_barrier_3_io_x_ppn;
  wire  tlb_entries_barrier_3_io_x_u;
  wire  tlb_entries_barrier_3_io_x_ae_ptw;
  wire  tlb_entries_barrier_3_io_x_ae_final;
  wire  tlb_entries_barrier_3_io_x_pf;
  wire  tlb_entries_barrier_3_io_x_gf;
  wire  tlb_entries_barrier_3_io_x_sw;
  wire  tlb_entries_barrier_3_io_x_sx;
  wire  tlb_entries_barrier_3_io_x_sr;
  wire  tlb_entries_barrier_3_io_x_pw;
  wire  tlb_entries_barrier_3_io_x_px;
  wire  tlb_entries_barrier_3_io_x_pr;
  wire  tlb_entries_barrier_3_io_x_ppp;
  wire  tlb_entries_barrier_3_io_x_pal;
  wire  tlb_entries_barrier_3_io_x_paa;
  wire  tlb_entries_barrier_3_io_x_eff;
  wire  tlb_entries_barrier_3_io_x_c;
  wire [19:0] tlb_entries_barrier_3_io_y_ppn;
  wire  tlb_entries_barrier_3_io_y_u;
  wire  tlb_entries_barrier_3_io_y_ae_ptw;
  wire  tlb_entries_barrier_3_io_y_ae_final;
  wire  tlb_entries_barrier_3_io_y_pf;
  wire  tlb_entries_barrier_3_io_y_gf;
  wire  tlb_entries_barrier_3_io_y_sw;
  wire  tlb_entries_barrier_3_io_y_sx;
  wire  tlb_entries_barrier_3_io_y_sr;
  wire  tlb_entries_barrier_3_io_y_pw;
  wire  tlb_entries_barrier_3_io_y_px;
  wire  tlb_entries_barrier_3_io_y_pr;
  wire  tlb_entries_barrier_3_io_y_ppp;
  wire  tlb_entries_barrier_3_io_y_pal;
  wire  tlb_entries_barrier_3_io_y_paa;
  wire  tlb_entries_barrier_3_io_y_eff;
  wire  tlb_entries_barrier_3_io_y_c;
  wire [19:0] tlb_entries_barrier_4_io_x_ppn;
  wire  tlb_entries_barrier_4_io_x_u;
  wire  tlb_entries_barrier_4_io_x_ae_ptw;
  wire  tlb_entries_barrier_4_io_x_ae_final;
  wire  tlb_entries_barrier_4_io_x_pf;
  wire  tlb_entries_barrier_4_io_x_gf;
  wire  tlb_entries_barrier_4_io_x_sw;
  wire  tlb_entries_barrier_4_io_x_sx;
  wire  tlb_entries_barrier_4_io_x_sr;
  wire  tlb_entries_barrier_4_io_x_pw;
  wire  tlb_entries_barrier_4_io_x_px;
  wire  tlb_entries_barrier_4_io_x_pr;
  wire  tlb_entries_barrier_4_io_x_ppp;
  wire  tlb_entries_barrier_4_io_x_pal;
  wire  tlb_entries_barrier_4_io_x_paa;
  wire  tlb_entries_barrier_4_io_x_eff;
  wire  tlb_entries_barrier_4_io_x_c;
  wire [19:0] tlb_entries_barrier_4_io_y_ppn;
  wire  tlb_entries_barrier_4_io_y_u;
  wire  tlb_entries_barrier_4_io_y_ae_ptw;
  wire  tlb_entries_barrier_4_io_y_ae_final;
  wire  tlb_entries_barrier_4_io_y_pf;
  wire  tlb_entries_barrier_4_io_y_gf;
  wire  tlb_entries_barrier_4_io_y_sw;
  wire  tlb_entries_barrier_4_io_y_sx;
  wire  tlb_entries_barrier_4_io_y_sr;
  wire  tlb_entries_barrier_4_io_y_pw;
  wire  tlb_entries_barrier_4_io_y_px;
  wire  tlb_entries_barrier_4_io_y_pr;
  wire  tlb_entries_barrier_4_io_y_ppp;
  wire  tlb_entries_barrier_4_io_y_pal;
  wire  tlb_entries_barrier_4_io_y_paa;
  wire  tlb_entries_barrier_4_io_y_eff;
  wire  tlb_entries_barrier_4_io_y_c;
  wire [19:0] tlb_entries_barrier_5_io_x_ppn;
  wire  tlb_entries_barrier_5_io_x_u;
  wire  tlb_entries_barrier_5_io_x_ae_ptw;
  wire  tlb_entries_barrier_5_io_x_ae_final;
  wire  tlb_entries_barrier_5_io_x_pf;
  wire  tlb_entries_barrier_5_io_x_gf;
  wire  tlb_entries_barrier_5_io_x_sw;
  wire  tlb_entries_barrier_5_io_x_sx;
  wire  tlb_entries_barrier_5_io_x_sr;
  wire  tlb_entries_barrier_5_io_x_pw;
  wire  tlb_entries_barrier_5_io_x_px;
  wire  tlb_entries_barrier_5_io_x_pr;
  wire  tlb_entries_barrier_5_io_x_ppp;
  wire  tlb_entries_barrier_5_io_x_pal;
  wire  tlb_entries_barrier_5_io_x_paa;
  wire  tlb_entries_barrier_5_io_x_eff;
  wire  tlb_entries_barrier_5_io_x_c;
  wire [19:0] tlb_entries_barrier_5_io_y_ppn;
  wire  tlb_entries_barrier_5_io_y_u;
  wire  tlb_entries_barrier_5_io_y_ae_ptw;
  wire  tlb_entries_barrier_5_io_y_ae_final;
  wire  tlb_entries_barrier_5_io_y_pf;
  wire  tlb_entries_barrier_5_io_y_gf;
  wire  tlb_entries_barrier_5_io_y_sw;
  wire  tlb_entries_barrier_5_io_y_sx;
  wire  tlb_entries_barrier_5_io_y_sr;
  wire  tlb_entries_barrier_5_io_y_pw;
  wire  tlb_entries_barrier_5_io_y_px;
  wire  tlb_entries_barrier_5_io_y_pr;
  wire  tlb_entries_barrier_5_io_y_ppp;
  wire  tlb_entries_barrier_5_io_y_pal;
  wire  tlb_entries_barrier_5_io_y_paa;
  wire  tlb_entries_barrier_5_io_y_eff;
  wire  tlb_entries_barrier_5_io_y_c;
  wire [19:0] tlb_entries_barrier_6_io_x_ppn;
  wire  tlb_entries_barrier_6_io_x_u;
  wire  tlb_entries_barrier_6_io_x_ae_ptw;
  wire  tlb_entries_barrier_6_io_x_ae_final;
  wire  tlb_entries_barrier_6_io_x_pf;
  wire  tlb_entries_barrier_6_io_x_gf;
  wire  tlb_entries_barrier_6_io_x_sw;
  wire  tlb_entries_barrier_6_io_x_sx;
  wire  tlb_entries_barrier_6_io_x_sr;
  wire  tlb_entries_barrier_6_io_x_pw;
  wire  tlb_entries_barrier_6_io_x_px;
  wire  tlb_entries_barrier_6_io_x_pr;
  wire  tlb_entries_barrier_6_io_x_ppp;
  wire  tlb_entries_barrier_6_io_x_pal;
  wire  tlb_entries_barrier_6_io_x_paa;
  wire  tlb_entries_barrier_6_io_x_eff;
  wire  tlb_entries_barrier_6_io_x_c;
  wire [19:0] tlb_entries_barrier_6_io_y_ppn;
  wire  tlb_entries_barrier_6_io_y_u;
  wire  tlb_entries_barrier_6_io_y_ae_ptw;
  wire  tlb_entries_barrier_6_io_y_ae_final;
  wire  tlb_entries_barrier_6_io_y_pf;
  wire  tlb_entries_barrier_6_io_y_gf;
  wire  tlb_entries_barrier_6_io_y_sw;
  wire  tlb_entries_barrier_6_io_y_sx;
  wire  tlb_entries_barrier_6_io_y_sr;
  wire  tlb_entries_barrier_6_io_y_pw;
  wire  tlb_entries_barrier_6_io_y_px;
  wire  tlb_entries_barrier_6_io_y_pr;
  wire  tlb_entries_barrier_6_io_y_ppp;
  wire  tlb_entries_barrier_6_io_y_pal;
  wire  tlb_entries_barrier_6_io_y_paa;
  wire  tlb_entries_barrier_6_io_y_eff;
  wire  tlb_entries_barrier_6_io_y_c;
  wire [19:0] tlb_entries_barrier_7_io_x_ppn;
  wire  tlb_entries_barrier_7_io_x_u;
  wire  tlb_entries_barrier_7_io_x_ae_ptw;
  wire  tlb_entries_barrier_7_io_x_ae_final;
  wire  tlb_entries_barrier_7_io_x_pf;
  wire  tlb_entries_barrier_7_io_x_gf;
  wire  tlb_entries_barrier_7_io_x_sw;
  wire  tlb_entries_barrier_7_io_x_sx;
  wire  tlb_entries_barrier_7_io_x_sr;
  wire  tlb_entries_barrier_7_io_x_pw;
  wire  tlb_entries_barrier_7_io_x_px;
  wire  tlb_entries_barrier_7_io_x_pr;
  wire  tlb_entries_barrier_7_io_x_ppp;
  wire  tlb_entries_barrier_7_io_x_pal;
  wire  tlb_entries_barrier_7_io_x_paa;
  wire  tlb_entries_barrier_7_io_x_eff;
  wire  tlb_entries_barrier_7_io_x_c;
  wire [19:0] tlb_entries_barrier_7_io_y_ppn;
  wire  tlb_entries_barrier_7_io_y_u;
  wire  tlb_entries_barrier_7_io_y_ae_ptw;
  wire  tlb_entries_barrier_7_io_y_ae_final;
  wire  tlb_entries_barrier_7_io_y_pf;
  wire  tlb_entries_barrier_7_io_y_gf;
  wire  tlb_entries_barrier_7_io_y_sw;
  wire  tlb_entries_barrier_7_io_y_sx;
  wire  tlb_entries_barrier_7_io_y_sr;
  wire  tlb_entries_barrier_7_io_y_pw;
  wire  tlb_entries_barrier_7_io_y_px;
  wire  tlb_entries_barrier_7_io_y_pr;
  wire  tlb_entries_barrier_7_io_y_ppp;
  wire  tlb_entries_barrier_7_io_y_pal;
  wire  tlb_entries_barrier_7_io_y_paa;
  wire  tlb_entries_barrier_7_io_y_eff;
  wire  tlb_entries_barrier_7_io_y_c;
  wire [19:0] tlb_entries_barrier_8_io_x_ppn;
  wire  tlb_entries_barrier_8_io_x_u;
  wire  tlb_entries_barrier_8_io_x_ae_ptw;
  wire  tlb_entries_barrier_8_io_x_ae_final;
  wire  tlb_entries_barrier_8_io_x_pf;
  wire  tlb_entries_barrier_8_io_x_gf;
  wire  tlb_entries_barrier_8_io_x_sw;
  wire  tlb_entries_barrier_8_io_x_sx;
  wire  tlb_entries_barrier_8_io_x_sr;
  wire  tlb_entries_barrier_8_io_x_pw;
  wire  tlb_entries_barrier_8_io_x_px;
  wire  tlb_entries_barrier_8_io_x_pr;
  wire  tlb_entries_barrier_8_io_x_ppp;
  wire  tlb_entries_barrier_8_io_x_pal;
  wire  tlb_entries_barrier_8_io_x_paa;
  wire  tlb_entries_barrier_8_io_x_eff;
  wire  tlb_entries_barrier_8_io_x_c;
  wire [19:0] tlb_entries_barrier_8_io_y_ppn;
  wire  tlb_entries_barrier_8_io_y_u;
  wire  tlb_entries_barrier_8_io_y_ae_ptw;
  wire  tlb_entries_barrier_8_io_y_ae_final;
  wire  tlb_entries_barrier_8_io_y_pf;
  wire  tlb_entries_barrier_8_io_y_gf;
  wire  tlb_entries_barrier_8_io_y_sw;
  wire  tlb_entries_barrier_8_io_y_sx;
  wire  tlb_entries_barrier_8_io_y_sr;
  wire  tlb_entries_barrier_8_io_y_pw;
  wire  tlb_entries_barrier_8_io_y_px;
  wire  tlb_entries_barrier_8_io_y_pr;
  wire  tlb_entries_barrier_8_io_y_ppp;
  wire  tlb_entries_barrier_8_io_y_pal;
  wire  tlb_entries_barrier_8_io_y_paa;
  wire  tlb_entries_barrier_8_io_y_eff;
  wire  tlb_entries_barrier_8_io_y_c;
  wire [19:0] tlb_entries_barrier_9_io_x_ppn;
  wire  tlb_entries_barrier_9_io_x_u;
  wire  tlb_entries_barrier_9_io_x_ae_ptw;
  wire  tlb_entries_barrier_9_io_x_ae_final;
  wire  tlb_entries_barrier_9_io_x_pf;
  wire  tlb_entries_barrier_9_io_x_gf;
  wire  tlb_entries_barrier_9_io_x_sw;
  wire  tlb_entries_barrier_9_io_x_sx;
  wire  tlb_entries_barrier_9_io_x_sr;
  wire  tlb_entries_barrier_9_io_x_pw;
  wire  tlb_entries_barrier_9_io_x_px;
  wire  tlb_entries_barrier_9_io_x_pr;
  wire  tlb_entries_barrier_9_io_x_ppp;
  wire  tlb_entries_barrier_9_io_x_pal;
  wire  tlb_entries_barrier_9_io_x_paa;
  wire  tlb_entries_barrier_9_io_x_eff;
  wire  tlb_entries_barrier_9_io_x_c;
  wire [19:0] tlb_entries_barrier_9_io_y_ppn;
  wire  tlb_entries_barrier_9_io_y_u;
  wire  tlb_entries_barrier_9_io_y_ae_ptw;
  wire  tlb_entries_barrier_9_io_y_ae_final;
  wire  tlb_entries_barrier_9_io_y_pf;
  wire  tlb_entries_barrier_9_io_y_gf;
  wire  tlb_entries_barrier_9_io_y_sw;
  wire  tlb_entries_barrier_9_io_y_sx;
  wire  tlb_entries_barrier_9_io_y_sr;
  wire  tlb_entries_barrier_9_io_y_pw;
  wire  tlb_entries_barrier_9_io_y_px;
  wire  tlb_entries_barrier_9_io_y_pr;
  wire  tlb_entries_barrier_9_io_y_ppp;
  wire  tlb_entries_barrier_9_io_y_pal;
  wire  tlb_entries_barrier_9_io_y_paa;
  wire  tlb_entries_barrier_9_io_y_eff;
  wire  tlb_entries_barrier_9_io_y_c;
  wire [19:0] tlb_entries_barrier_10_io_x_ppn;
  wire  tlb_entries_barrier_10_io_x_u;
  wire  tlb_entries_barrier_10_io_x_ae_ptw;
  wire  tlb_entries_barrier_10_io_x_ae_final;
  wire  tlb_entries_barrier_10_io_x_pf;
  wire  tlb_entries_barrier_10_io_x_gf;
  wire  tlb_entries_barrier_10_io_x_sw;
  wire  tlb_entries_barrier_10_io_x_sx;
  wire  tlb_entries_barrier_10_io_x_sr;
  wire  tlb_entries_barrier_10_io_x_pw;
  wire  tlb_entries_barrier_10_io_x_px;
  wire  tlb_entries_barrier_10_io_x_pr;
  wire  tlb_entries_barrier_10_io_x_ppp;
  wire  tlb_entries_barrier_10_io_x_pal;
  wire  tlb_entries_barrier_10_io_x_paa;
  wire  tlb_entries_barrier_10_io_x_eff;
  wire  tlb_entries_barrier_10_io_x_c;
  wire [19:0] tlb_entries_barrier_10_io_y_ppn;
  wire  tlb_entries_barrier_10_io_y_u;
  wire  tlb_entries_barrier_10_io_y_ae_ptw;
  wire  tlb_entries_barrier_10_io_y_ae_final;
  wire  tlb_entries_barrier_10_io_y_pf;
  wire  tlb_entries_barrier_10_io_y_gf;
  wire  tlb_entries_barrier_10_io_y_sw;
  wire  tlb_entries_barrier_10_io_y_sx;
  wire  tlb_entries_barrier_10_io_y_sr;
  wire  tlb_entries_barrier_10_io_y_pw;
  wire  tlb_entries_barrier_10_io_y_px;
  wire  tlb_entries_barrier_10_io_y_pr;
  wire  tlb_entries_barrier_10_io_y_ppp;
  wire  tlb_entries_barrier_10_io_y_pal;
  wire  tlb_entries_barrier_10_io_y_paa;
  wire  tlb_entries_barrier_10_io_y_eff;
  wire  tlb_entries_barrier_10_io_y_c;
  wire [19:0] tlb_entries_barrier_11_io_x_ppn;
  wire  tlb_entries_barrier_11_io_x_u;
  wire  tlb_entries_barrier_11_io_x_ae_ptw;
  wire  tlb_entries_barrier_11_io_x_ae_final;
  wire  tlb_entries_barrier_11_io_x_pf;
  wire  tlb_entries_barrier_11_io_x_gf;
  wire  tlb_entries_barrier_11_io_x_sw;
  wire  tlb_entries_barrier_11_io_x_sx;
  wire  tlb_entries_barrier_11_io_x_sr;
  wire  tlb_entries_barrier_11_io_x_pw;
  wire  tlb_entries_barrier_11_io_x_px;
  wire  tlb_entries_barrier_11_io_x_pr;
  wire  tlb_entries_barrier_11_io_x_ppp;
  wire  tlb_entries_barrier_11_io_x_pal;
  wire  tlb_entries_barrier_11_io_x_paa;
  wire  tlb_entries_barrier_11_io_x_eff;
  wire  tlb_entries_barrier_11_io_x_c;
  wire [19:0] tlb_entries_barrier_11_io_y_ppn;
  wire  tlb_entries_barrier_11_io_y_u;
  wire  tlb_entries_barrier_11_io_y_ae_ptw;
  wire  tlb_entries_barrier_11_io_y_ae_final;
  wire  tlb_entries_barrier_11_io_y_pf;
  wire  tlb_entries_barrier_11_io_y_gf;
  wire  tlb_entries_barrier_11_io_y_sw;
  wire  tlb_entries_barrier_11_io_y_sx;
  wire  tlb_entries_barrier_11_io_y_sr;
  wire  tlb_entries_barrier_11_io_y_pw;
  wire  tlb_entries_barrier_11_io_y_px;
  wire  tlb_entries_barrier_11_io_y_pr;
  wire  tlb_entries_barrier_11_io_y_ppp;
  wire  tlb_entries_barrier_11_io_y_pal;
  wire  tlb_entries_barrier_11_io_y_paa;
  wire  tlb_entries_barrier_11_io_y_eff;
  wire  tlb_entries_barrier_11_io_y_c;
  wire [19:0] tlb_entries_barrier_12_io_x_ppn;
  wire  tlb_entries_barrier_12_io_x_u;
  wire  tlb_entries_barrier_12_io_x_ae_ptw;
  wire  tlb_entries_barrier_12_io_x_ae_final;
  wire  tlb_entries_barrier_12_io_x_pf;
  wire  tlb_entries_barrier_12_io_x_gf;
  wire  tlb_entries_barrier_12_io_x_sw;
  wire  tlb_entries_barrier_12_io_x_sx;
  wire  tlb_entries_barrier_12_io_x_sr;
  wire  tlb_entries_barrier_12_io_x_pw;
  wire  tlb_entries_barrier_12_io_x_px;
  wire  tlb_entries_barrier_12_io_x_pr;
  wire  tlb_entries_barrier_12_io_x_ppp;
  wire  tlb_entries_barrier_12_io_x_pal;
  wire  tlb_entries_barrier_12_io_x_paa;
  wire  tlb_entries_barrier_12_io_x_eff;
  wire  tlb_entries_barrier_12_io_x_c;
  wire [19:0] tlb_entries_barrier_12_io_y_ppn;
  wire  tlb_entries_barrier_12_io_y_u;
  wire  tlb_entries_barrier_12_io_y_ae_ptw;
  wire  tlb_entries_barrier_12_io_y_ae_final;
  wire  tlb_entries_barrier_12_io_y_pf;
  wire  tlb_entries_barrier_12_io_y_gf;
  wire  tlb_entries_barrier_12_io_y_sw;
  wire  tlb_entries_barrier_12_io_y_sx;
  wire  tlb_entries_barrier_12_io_y_sr;
  wire  tlb_entries_barrier_12_io_y_pw;
  wire  tlb_entries_barrier_12_io_y_px;
  wire  tlb_entries_barrier_12_io_y_pr;
  wire  tlb_entries_barrier_12_io_y_ppp;
  wire  tlb_entries_barrier_12_io_y_pal;
  wire  tlb_entries_barrier_12_io_y_paa;
  wire  tlb_entries_barrier_12_io_y_eff;
  wire  tlb_entries_barrier_12_io_y_c;
  wire [19:0] tlb_vpn = tlb_io_req_bits_vaddr[31:12];
  reg [19:0] tlb_sectored_entries_0_0_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_0_data_0;
  reg [40:0] tlb_sectored_entries_0_0_data_1;
  reg [40:0] tlb_sectored_entries_0_0_data_2;
  reg [40:0] tlb_sectored_entries_0_0_data_3;
  reg  tlb_sectored_entries_0_0_valid_0;
  reg  tlb_sectored_entries_0_0_valid_1;
  reg  tlb_sectored_entries_0_0_valid_2;
  reg  tlb_sectored_entries_0_0_valid_3;
  reg [19:0] tlb_sectored_entries_0_1_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_1_data_0;
  reg [40:0] tlb_sectored_entries_0_1_data_1;
  reg [40:0] tlb_sectored_entries_0_1_data_2;
  reg [40:0] tlb_sectored_entries_0_1_data_3;
  reg  tlb_sectored_entries_0_1_valid_0;
  reg  tlb_sectored_entries_0_1_valid_1;
  reg  tlb_sectored_entries_0_1_valid_2;
  reg  tlb_sectored_entries_0_1_valid_3;
  reg [19:0] tlb_sectored_entries_0_2_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_2_data_0;
  reg [40:0] tlb_sectored_entries_0_2_data_1;
  reg [40:0] tlb_sectored_entries_0_2_data_2;
  reg [40:0] tlb_sectored_entries_0_2_data_3;
  reg  tlb_sectored_entries_0_2_valid_0;
  reg  tlb_sectored_entries_0_2_valid_1;
  reg  tlb_sectored_entries_0_2_valid_2;
  reg  tlb_sectored_entries_0_2_valid_3;
  reg [19:0] tlb_sectored_entries_0_3_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_3_data_0;
  reg [40:0] tlb_sectored_entries_0_3_data_1;
  reg [40:0] tlb_sectored_entries_0_3_data_2;
  reg [40:0] tlb_sectored_entries_0_3_data_3;
  reg  tlb_sectored_entries_0_3_valid_0;
  reg  tlb_sectored_entries_0_3_valid_1;
  reg  tlb_sectored_entries_0_3_valid_2;
  reg  tlb_sectored_entries_0_3_valid_3;
  reg [19:0] tlb_sectored_entries_0_4_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_4_data_0;
  reg [40:0] tlb_sectored_entries_0_4_data_1;
  reg [40:0] tlb_sectored_entries_0_4_data_2;
  reg [40:0] tlb_sectored_entries_0_4_data_3;
  reg  tlb_sectored_entries_0_4_valid_0;
  reg  tlb_sectored_entries_0_4_valid_1;
  reg  tlb_sectored_entries_0_4_valid_2;
  reg  tlb_sectored_entries_0_4_valid_3;
  reg [19:0] tlb_sectored_entries_0_5_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_5_data_0;
  reg [40:0] tlb_sectored_entries_0_5_data_1;
  reg [40:0] tlb_sectored_entries_0_5_data_2;
  reg [40:0] tlb_sectored_entries_0_5_data_3;
  reg  tlb_sectored_entries_0_5_valid_0;
  reg  tlb_sectored_entries_0_5_valid_1;
  reg  tlb_sectored_entries_0_5_valid_2;
  reg  tlb_sectored_entries_0_5_valid_3;
  reg [19:0] tlb_sectored_entries_0_6_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_6_data_0;
  reg [40:0] tlb_sectored_entries_0_6_data_1;
  reg [40:0] tlb_sectored_entries_0_6_data_2;
  reg [40:0] tlb_sectored_entries_0_6_data_3;
  reg  tlb_sectored_entries_0_6_valid_0;
  reg  tlb_sectored_entries_0_6_valid_1;
  reg  tlb_sectored_entries_0_6_valid_2;
  reg  tlb_sectored_entries_0_6_valid_3;
  reg [19:0] tlb_sectored_entries_0_7_tag_vpn;
  reg [40:0] tlb_sectored_entries_0_7_data_0;
  reg [40:0] tlb_sectored_entries_0_7_data_1;
  reg [40:0] tlb_sectored_entries_0_7_data_2;
  reg [40:0] tlb_sectored_entries_0_7_data_3;
  reg  tlb_sectored_entries_0_7_valid_0;
  reg  tlb_sectored_entries_0_7_valid_1;
  reg  tlb_sectored_entries_0_7_valid_2;
  reg  tlb_sectored_entries_0_7_valid_3;
  reg [19:0] tlb_superpage_entries_0_tag_vpn;
  reg [40:0] tlb_superpage_entries_0_data_0;
  reg  tlb_superpage_entries_0_valid_0;
  reg [19:0] tlb_superpage_entries_1_tag_vpn;
  reg [40:0] tlb_superpage_entries_1_data_0;
  reg  tlb_superpage_entries_1_valid_0;
  reg [19:0] tlb_superpage_entries_2_tag_vpn;
  reg [40:0] tlb_superpage_entries_2_data_0;
  reg  tlb_superpage_entries_2_valid_0;
  reg [19:0] tlb_superpage_entries_3_tag_vpn;
  reg [40:0] tlb_superpage_entries_3_data_0;
  reg  tlb_superpage_entries_3_valid_0;
  reg  tlb_special_entry_level;
  reg [19:0] tlb_special_entry_tag_vpn;
  reg [40:0] tlb_special_entry_data_0;
  reg  tlb_special_entry_valid_0;
  reg [1:0] tlb_state;
  reg [19:0] tlb_r_refill_tag;
  reg [1:0] tlb_r_superpage_repl_addr;
  reg [2:0] tlb_r_sectored_repl_addr;
  reg  tlb_r_sectored_hit_valid;
  reg [2:0] tlb_r_sectored_hit_bits;
  reg  tlb_r_need_gpa;
  wire  tlb_priv_s = tlb_io_req_bits_prv[0];
  wire  tlb_priv_uses_vm = tlb_io_req_bits_prv <= 2'h1;
  wire  tlb__vm_enabled_T_1 = tlb_io_ptw_ptbr_mode & tlb_priv_uses_vm;
  wire  tlb__vm_enabled_T_2 = ~tlb_io_req_bits_passthrough;
  wire  tlb_vm_enabled = tlb__vm_enabled_T_1 & tlb__vm_enabled_T_2;
  wire [19:0] tlb_refill_ppn = tlb_io_ptw_resp_bits_pte_ppn[19:0];
  wire  tlb__invalidate_refill_T = tlb_state == 2'h1;
  wire  tlb__invalidate_refill_T_1 = tlb_state == 2'h3;
  wire  tlb__invalidate_refill_T_2 = tlb__invalidate_refill_T | tlb__invalidate_refill_T_1;
  wire  tlb_invalidate_refill = tlb__invalidate_refill_T_2 | tlb_io_sfence_valid;
  wire  tlb__mpu_ppn_T_20 = tlb_special_entry_data_0[19];
  wire [9:0] tlb_mpu_ppn_res = tlb_mpu_ppn_barrier_io_y_ppn[19:10];
  wire  tlb__mpu_ppn_ignore_T = tlb_special_entry_level < 1'h1;
  wire [19:0] tlb__mpu_ppn_T_23 = tlb__mpu_ppn_ignore_T ? tlb_vpn : 20'h0;
  wire [19:0] tlb__mpu_ppn_T_24 = tlb__mpu_ppn_T_23 | tlb_mpu_ppn_barrier_io_y_ppn;
  wire [9:0] tlb__mpu_ppn_T_25 = tlb__mpu_ppn_T_24[9:0];
  wire [19:0] tlb__mpu_ppn_T_26 = {tlb_mpu_ppn_res,tlb__mpu_ppn_T_25};
  wire [19:0] tlb__mpu_ppn_T_27 = tlb_io_req_bits_vaddr[31:12];
  wire [19:0] tlb__mpu_ppn_T_28 = tlb_vm_enabled ? tlb__mpu_ppn_T_26 : tlb__mpu_ppn_T_27;
  wire [19:0] tlb_mpu_ppn = tlb_io_ptw_resp_valid ? tlb_refill_ppn : tlb__mpu_ppn_T_28;
  wire [11:0] tlb__mpu_physaddr_T = tlb_io_req_bits_vaddr[11:0];
  wire [31:0] tlb_mpu_physaddr = {tlb_mpu_ppn,tlb__mpu_physaddr_T};
  wire  tlb__mpu_priv_T = tlb_io_ptw_resp_valid | tlb_io_req_bits_passthrough;
  wire [2:0] tlb__mpu_priv_T_2 = {tlb_io_ptw_status_debug,tlb_io_req_bits_prv};
  wire [2:0] tlb_mpu_priv = tlb__mpu_priv_T ? 3'h1 : tlb__mpu_priv_T_2;
  wire [31:0] tlb__legal_address_T = tlb_mpu_physaddr ^ 32'h3000;
  wire [32:0] tlb__legal_address_T_1 = {1'b0,$signed(tlb__legal_address_T)};
  wire [32:0] tlb__legal_address_T_3 = $signed(tlb__legal_address_T_1) & -33'sh1000;
  wire  tlb__legal_address_T_4 = $signed(tlb__legal_address_T_3) == 33'sh0;
  wire [31:0] tlb__legal_address_T_5 = tlb_mpu_physaddr ^ 32'hc000000;
  wire [32:0] tlb__legal_address_T_6 = {1'b0,$signed(tlb__legal_address_T_5)};
  wire [32:0] tlb__legal_address_T_8 = $signed(tlb__legal_address_T_6) & -33'sh4000000;
  wire  tlb__legal_address_T_9 = $signed(tlb__legal_address_T_8) == 33'sh0;
  wire [31:0] tlb__legal_address_T_10 = tlb_mpu_physaddr ^ 32'h2000000;
  wire [32:0] tlb__legal_address_T_11 = {1'b0,$signed(tlb__legal_address_T_10)};
  wire [32:0] tlb__legal_address_T_13 = $signed(tlb__legal_address_T_11) & -33'sh10000;
  wire  tlb__legal_address_T_14 = $signed(tlb__legal_address_T_13) == 33'sh0;
  wire [32:0] tlb__legal_address_T_16 = {1'b0,$signed(tlb_mpu_physaddr)};
  wire [32:0] tlb__legal_address_T_18 = $signed(tlb__legal_address_T_16) & -33'sh1000;
  wire  tlb__legal_address_T_19 = $signed(tlb__legal_address_T_18) == 33'sh0;
  wire [31:0] tlb__legal_address_T_20 = tlb_mpu_physaddr ^ 32'h10000;
  wire [32:0] tlb__legal_address_T_21 = {1'b0,$signed(tlb__legal_address_T_20)};
  wire [32:0] tlb__legal_address_T_23 = $signed(tlb__legal_address_T_21) & -33'sh10000;
  wire  tlb__legal_address_T_24 = $signed(tlb__legal_address_T_23) == 33'sh0;
  wire [31:0] tlb__legal_address_T_25 = tlb_mpu_physaddr ^ 32'h10000000;
  wire [32:0] tlb__legal_address_T_26 = {1'b0,$signed(tlb__legal_address_T_25)};
  wire [32:0] tlb__legal_address_T_28 = $signed(tlb__legal_address_T_26) & -33'sh10000000;
  wire  tlb__legal_address_T_29 = $signed(tlb__legal_address_T_28) == 33'sh0;
  wire [31:0] tlb__legal_address_T_30 = tlb_mpu_physaddr ^ 32'h20000000;
  wire [32:0] tlb__legal_address_T_31 = {1'b0,$signed(tlb__legal_address_T_30)};
  wire [32:0] tlb__legal_address_T_33 = $signed(tlb__legal_address_T_31) & -33'sh20000000;
  wire  tlb__legal_address_T_34 = $signed(tlb__legal_address_T_33) == 33'sh0;
  wire [31:0] tlb__legal_address_T_35 = tlb_mpu_physaddr ^ 32'h40000000;
  wire [32:0] tlb__legal_address_T_36 = {1'b0,$signed(tlb__legal_address_T_35)};
  wire [32:0] tlb__legal_address_T_38 = $signed(tlb__legal_address_T_36) & -33'sh40000000;
  wire  tlb__legal_address_T_39 = $signed(tlb__legal_address_T_38) == 33'sh0;
  wire [31:0] tlb__legal_address_T_40 = tlb_mpu_physaddr ^ 32'h80000000;
  wire [32:0] tlb__legal_address_T_41 = {1'b0,$signed(tlb__legal_address_T_40)};
  wire [32:0] tlb__legal_address_T_43 = $signed(tlb__legal_address_T_41) & -33'sh40000000;
  wire  tlb__legal_address_T_44 = $signed(tlb__legal_address_T_43) == 33'sh0;
  wire  tlb__legal_address_T_45 = tlb__legal_address_T_29 | tlb__legal_address_T_34;
  wire  tlb__legal_address_T_46 = tlb__legal_address_T_45 | tlb__legal_address_T_39;
  wire  tlb__legal_address_T_47 = tlb__legal_address_T_46 | tlb__legal_address_T_44;
  wire [31:0] tlb__legal_address_T_48 = tlb_mpu_physaddr ^ 32'hc0000000;
  wire [32:0] tlb__legal_address_T_49 = {1'b0,$signed(tlb__legal_address_T_48)};
  wire [32:0] tlb__legal_address_T_51 = $signed(tlb__legal_address_T_49) & -33'sh40000000;
  wire  tlb__legal_address_T_52 = $signed(tlb__legal_address_T_51) == 33'sh0;
  wire  tlb__legal_address_T_53 = tlb__legal_address_T_4 | tlb__legal_address_T_9;
  wire  tlb__legal_address_T_54 = tlb__legal_address_T_53 | tlb__legal_address_T_14;
  wire  tlb__legal_address_T_55 = tlb__legal_address_T_54 | tlb__legal_address_T_19;
  wire  tlb__legal_address_T_56 = tlb__legal_address_T_55 | tlb__legal_address_T_24;
  wire  tlb__legal_address_T_57 = tlb__legal_address_T_56 | tlb__legal_address_T_47;
  wire  tlb_legal_address = tlb__legal_address_T_57 | tlb__legal_address_T_52;
  wire [32:0] tlb__cacheable_T_3 = $signed(tlb__legal_address_T_16) & 33'shf8010000;
  wire  tlb__cacheable_T_4 = $signed(tlb__cacheable_T_3) == 33'sh0;
  wire [31:0] tlb__cacheable_T_5 = tlb_mpu_physaddr ^ 32'h8000000;
  wire [32:0] tlb__cacheable_T_6 = {1'b0,$signed(tlb__cacheable_T_5)};
  wire [32:0] tlb__cacheable_T_8 = $signed(tlb__cacheable_T_6) & 33'shf8000000;
  wire  tlb__cacheable_T_9 = $signed(tlb__cacheable_T_8) == 33'sh0;
  wire [32:0] tlb__cacheable_T_13 = $signed(tlb__legal_address_T_49) & 33'shc0000000;
  wire  tlb__cacheable_T_14 = $signed(tlb__cacheable_T_13) == 33'sh0;
  wire  tlb__cacheable_T_15 = tlb__cacheable_T_4 | tlb__cacheable_T_9;
  wire [32:0] tlb__cacheable_T_20 = $signed(tlb__legal_address_T_21) & 33'shf8010000;
  wire  tlb__cacheable_T_21 = $signed(tlb__cacheable_T_20) == 33'sh0;
  wire [32:0] tlb__cacheable_T_25 = $signed(tlb__legal_address_T_26) & 33'shf0000000;
  wire  tlb__cacheable_T_26 = $signed(tlb__cacheable_T_25) == 33'sh0;
  wire [32:0] tlb__cacheable_T_30 = $signed(tlb__legal_address_T_31) & 33'she0000000;
  wire  tlb__cacheable_T_31 = $signed(tlb__cacheable_T_30) == 33'sh0;
  wire [32:0] tlb__cacheable_T_35 = $signed(tlb__legal_address_T_36) & 33'shc0000000;
  wire  tlb__cacheable_T_36 = $signed(tlb__cacheable_T_35) == 33'sh0;
  wire [32:0] tlb__cacheable_T_40 = $signed(tlb__legal_address_T_41) & 33'shc0000000;
  wire  tlb__cacheable_T_41 = $signed(tlb__cacheable_T_40) == 33'sh0;
  wire  tlb__cacheable_T_42 = tlb__cacheable_T_21 | tlb__cacheable_T_26;
  wire  tlb__cacheable_T_43 = tlb__cacheable_T_42 | tlb__cacheable_T_31;
  wire  tlb__cacheable_T_44 = tlb__cacheable_T_43 | tlb__cacheable_T_36;
  wire  tlb__cacheable_T_45 = tlb__cacheable_T_44 | tlb__cacheable_T_41;
  wire  tlb__cacheable_T_49 = tlb_legal_address & tlb__cacheable_T_45;
  wire  tlb__deny_access_to_debug_T = tlb_mpu_priv <= 3'h3;
  wire  tlb_deny_access_to_debug = tlb__deny_access_to_debug_T & tlb__legal_address_T_19;
  wire  tlb__prot_r_T_6 = ~tlb_deny_access_to_debug;
  wire  tlb__prot_r_T_7 = tlb_legal_address & tlb__prot_r_T_6;
  wire  tlb_prot_r = tlb__prot_r_T_7 & tlb_pmp_io_r;
  wire [32:0] tlb__prot_w_T_28 = $signed(tlb__legal_address_T_41) & 33'sh80000000;
  wire  tlb__prot_w_T_29 = $signed(tlb__prot_w_T_28) == 33'sh0;
  wire  tlb__prot_w_T_31 = tlb__cacheable_T_15 | tlb__cacheable_T_26;
  wire  tlb__prot_w_T_32 = tlb__prot_w_T_31 | tlb__cacheable_T_31;
  wire  tlb__prot_w_T_33 = tlb__prot_w_T_32 | tlb__cacheable_T_36;
  wire  tlb__prot_w_T_34 = tlb__prot_w_T_33 | tlb__prot_w_T_29;
  wire  tlb__prot_w_T_43 = tlb_legal_address & tlb__prot_w_T_34;
  wire  tlb__prot_w_T_45 = tlb__prot_w_T_43 & tlb__prot_r_T_6;
  wire  tlb_prot_w = tlb__prot_w_T_45 & tlb_pmp_io_w;
  wire  tlb_prot_al = tlb_legal_address & tlb__cacheable_T_15;
  wire [32:0] tlb__prot_x_T_3 = $signed(tlb__legal_address_T_16) & 33'shfa000000;
  wire  tlb__prot_x_T_4 = $signed(tlb__prot_x_T_3) == 33'sh0;
  wire  tlb__prot_x_T_25 = tlb__prot_x_T_4 | tlb__cacheable_T_26;
  wire  tlb__prot_x_T_26 = tlb__prot_x_T_25 | tlb__cacheable_T_31;
  wire  tlb__prot_x_T_27 = tlb__prot_x_T_26 | tlb__cacheable_T_36;
  wire  tlb__prot_x_T_28 = tlb__prot_x_T_27 | tlb__prot_w_T_29;
  wire  tlb__prot_x_T_43 = tlb_legal_address & tlb__prot_x_T_28;
  wire  tlb__prot_x_T_45 = tlb__prot_x_T_43 & tlb__prot_r_T_6;
  wire  tlb_prot_x = tlb__prot_x_T_45 & tlb_pmp_io_x;
  wire [32:0] tlb__prot_eff_T_38 = $signed(tlb__legal_address_T_16) & 33'shfa012000;
  wire  tlb__prot_eff_T_39 = $signed(tlb__prot_eff_T_38) == 33'sh0;
  wire [32:0] tlb__prot_eff_T_43 = $signed(tlb__legal_address_T_11) & 33'shfa010000;
  wire  tlb__prot_eff_T_44 = $signed(tlb__prot_eff_T_43) == 33'sh0;
  wire  tlb__prot_eff_T_55 = tlb__prot_eff_T_39 | tlb__prot_eff_T_44;
  wire  tlb__prot_eff_T_56 = tlb__prot_eff_T_55 | tlb__cacheable_T_9;
  wire  tlb__prot_eff_T_57 = tlb__prot_eff_T_56 | tlb__cacheable_T_14;
  wire  tlb_prot_eff = tlb_legal_address & tlb__prot_eff_T_57;
  wire  tlb__sector_hits_T = tlb_sectored_entries_0_0_valid_0 | tlb_sectored_entries_0_0_valid_1;
  wire  tlb__sector_hits_T_1 = tlb__sector_hits_T | tlb_sectored_entries_0_0_valid_2;
  wire  tlb__sector_hits_T_2 = tlb__sector_hits_T_1 | tlb_sectored_entries_0_0_valid_3;
  wire [19:0] tlb__sector_hits_T_3 = tlb_sectored_entries_0_0_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_4 = tlb__sector_hits_T_3[19:2];
  wire  tlb__sector_hits_T_5 = tlb__sector_hits_T_4 == 18'h0;
  wire  tlb_sector_hits_0 = tlb__sector_hits_T_2 & tlb__sector_hits_T_5;
  wire  tlb__sector_hits_T_8 = tlb_sectored_entries_0_1_valid_0 | tlb_sectored_entries_0_1_valid_1;
  wire  tlb__sector_hits_T_9 = tlb__sector_hits_T_8 | tlb_sectored_entries_0_1_valid_2;
  wire  tlb__sector_hits_T_10 = tlb__sector_hits_T_9 | tlb_sectored_entries_0_1_valid_3;
  wire [19:0] tlb__sector_hits_T_11 = tlb_sectored_entries_0_1_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_12 = tlb__sector_hits_T_11[19:2];
  wire  tlb__sector_hits_T_13 = tlb__sector_hits_T_12 == 18'h0;
  wire  tlb_sector_hits_1 = tlb__sector_hits_T_10 & tlb__sector_hits_T_13;
  wire  tlb__sector_hits_T_16 = tlb_sectored_entries_0_2_valid_0 | tlb_sectored_entries_0_2_valid_1;
  wire  tlb__sector_hits_T_17 = tlb__sector_hits_T_16 | tlb_sectored_entries_0_2_valid_2;
  wire  tlb__sector_hits_T_18 = tlb__sector_hits_T_17 | tlb_sectored_entries_0_2_valid_3;
  wire [19:0] tlb__sector_hits_T_19 = tlb_sectored_entries_0_2_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_20 = tlb__sector_hits_T_19[19:2];
  wire  tlb__sector_hits_T_21 = tlb__sector_hits_T_20 == 18'h0;
  wire  tlb_sector_hits_2 = tlb__sector_hits_T_18 & tlb__sector_hits_T_21;
  wire  tlb__sector_hits_T_24 = tlb_sectored_entries_0_3_valid_0 | tlb_sectored_entries_0_3_valid_1;
  wire  tlb__sector_hits_T_25 = tlb__sector_hits_T_24 | tlb_sectored_entries_0_3_valid_2;
  wire  tlb__sector_hits_T_26 = tlb__sector_hits_T_25 | tlb_sectored_entries_0_3_valid_3;
  wire [19:0] tlb__sector_hits_T_27 = tlb_sectored_entries_0_3_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_28 = tlb__sector_hits_T_27[19:2];
  wire  tlb__sector_hits_T_29 = tlb__sector_hits_T_28 == 18'h0;
  wire  tlb_sector_hits_3 = tlb__sector_hits_T_26 & tlb__sector_hits_T_29;
  wire  tlb__sector_hits_T_32 = tlb_sectored_entries_0_4_valid_0 | tlb_sectored_entries_0_4_valid_1;
  wire  tlb__sector_hits_T_33 = tlb__sector_hits_T_32 | tlb_sectored_entries_0_4_valid_2;
  wire  tlb__sector_hits_T_34 = tlb__sector_hits_T_33 | tlb_sectored_entries_0_4_valid_3;
  wire [19:0] tlb__sector_hits_T_35 = tlb_sectored_entries_0_4_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_36 = tlb__sector_hits_T_35[19:2];
  wire  tlb__sector_hits_T_37 = tlb__sector_hits_T_36 == 18'h0;
  wire  tlb_sector_hits_4 = tlb__sector_hits_T_34 & tlb__sector_hits_T_37;
  wire  tlb__sector_hits_T_40 = tlb_sectored_entries_0_5_valid_0 | tlb_sectored_entries_0_5_valid_1;
  wire  tlb__sector_hits_T_41 = tlb__sector_hits_T_40 | tlb_sectored_entries_0_5_valid_2;
  wire  tlb__sector_hits_T_42 = tlb__sector_hits_T_41 | tlb_sectored_entries_0_5_valid_3;
  wire [19:0] tlb__sector_hits_T_43 = tlb_sectored_entries_0_5_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_44 = tlb__sector_hits_T_43[19:2];
  wire  tlb__sector_hits_T_45 = tlb__sector_hits_T_44 == 18'h0;
  wire  tlb_sector_hits_5 = tlb__sector_hits_T_42 & tlb__sector_hits_T_45;
  wire  tlb__sector_hits_T_48 = tlb_sectored_entries_0_6_valid_0 | tlb_sectored_entries_0_6_valid_1;
  wire  tlb__sector_hits_T_49 = tlb__sector_hits_T_48 | tlb_sectored_entries_0_6_valid_2;
  wire  tlb__sector_hits_T_50 = tlb__sector_hits_T_49 | tlb_sectored_entries_0_6_valid_3;
  wire [19:0] tlb__sector_hits_T_51 = tlb_sectored_entries_0_6_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_52 = tlb__sector_hits_T_51[19:2];
  wire  tlb__sector_hits_T_53 = tlb__sector_hits_T_52 == 18'h0;
  wire  tlb_sector_hits_6 = tlb__sector_hits_T_50 & tlb__sector_hits_T_53;
  wire  tlb__sector_hits_T_56 = tlb_sectored_entries_0_7_valid_0 | tlb_sectored_entries_0_7_valid_1;
  wire  tlb__sector_hits_T_57 = tlb__sector_hits_T_56 | tlb_sectored_entries_0_7_valid_2;
  wire  tlb__sector_hits_T_58 = tlb__sector_hits_T_57 | tlb_sectored_entries_0_7_valid_3;
  wire [19:0] tlb__sector_hits_T_59 = tlb_sectored_entries_0_7_tag_vpn ^ tlb_vpn;
  wire [17:0] tlb__sector_hits_T_60 = tlb__sector_hits_T_59[19:2];
  wire  tlb__sector_hits_T_61 = tlb__sector_hits_T_60 == 18'h0;
  wire  tlb_sector_hits_7 = tlb__sector_hits_T_58 & tlb__sector_hits_T_61;
  wire [19:0] tlb__superpage_hits_T = tlb_superpage_entries_0_tag_vpn ^ tlb_vpn;
  wire [9:0] tlb__superpage_hits_T_1 = tlb__superpage_hits_T[19:10];
  wire  tlb__superpage_hits_T_2 = tlb__superpage_hits_T_1 == 10'h0;
  wire  tlb__superpage_hits_T_4 = tlb_superpage_entries_0_valid_0 & tlb__superpage_hits_T_2;
  wire [19:0] tlb__superpage_hits_T_9 = tlb_superpage_entries_1_tag_vpn ^ tlb_vpn;
  wire [9:0] tlb__superpage_hits_T_10 = tlb__superpage_hits_T_9[19:10];
  wire  tlb__superpage_hits_T_11 = tlb__superpage_hits_T_10 == 10'h0;
  wire  tlb__superpage_hits_T_13 = tlb_superpage_entries_1_valid_0 & tlb__superpage_hits_T_11;
  wire [19:0] tlb__superpage_hits_T_18 = tlb_superpage_entries_2_tag_vpn ^ tlb_vpn;
  wire [9:0] tlb__superpage_hits_T_19 = tlb__superpage_hits_T_18[19:10];
  wire  tlb__superpage_hits_T_20 = tlb__superpage_hits_T_19 == 10'h0;
  wire  tlb__superpage_hits_T_22 = tlb_superpage_entries_2_valid_0 & tlb__superpage_hits_T_20;
  wire [19:0] tlb__superpage_hits_T_27 = tlb_superpage_entries_3_tag_vpn ^ tlb_vpn;
  wire [9:0] tlb__superpage_hits_T_28 = tlb__superpage_hits_T_27[19:10];
  wire  tlb__superpage_hits_T_29 = tlb__superpage_hits_T_28 == 10'h0;
  wire  tlb__superpage_hits_T_31 = tlb_superpage_entries_3_valid_0 & tlb__superpage_hits_T_29;
  wire [1:0] tlb_hitsVec_idx = tlb_vpn[1:0];
  wire  tlb__GEN_1 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_0_valid_1 : tlb_sectored_entries_0_0_valid_0;
  wire  tlb__GEN_2 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_0_valid_2 : tlb__GEN_1;
  wire  tlb__GEN_3 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_0_valid_3 : tlb__GEN_2;
  wire  tlb__hitsVec_T_5 = tlb__GEN_3 & tlb__sector_hits_T_5;
  wire  tlb_hitsVec_0 = tlb_vm_enabled & tlb__hitsVec_T_5;
  wire  tlb__GEN_5 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_1_valid_1 : tlb_sectored_entries_0_1_valid_0;
  wire  tlb__GEN_6 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_1_valid_2 : tlb__GEN_5;
  wire  tlb__GEN_7 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_1_valid_3 : tlb__GEN_6;
  wire  tlb__hitsVec_T_11 = tlb__GEN_7 & tlb__sector_hits_T_13;
  wire  tlb_hitsVec_1 = tlb_vm_enabled & tlb__hitsVec_T_11;
  wire  tlb__GEN_9 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_2_valid_1 : tlb_sectored_entries_0_2_valid_0;
  wire  tlb__GEN_10 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_2_valid_2 : tlb__GEN_9;
  wire  tlb__GEN_11 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_2_valid_3 : tlb__GEN_10;
  wire  tlb__hitsVec_T_17 = tlb__GEN_11 & tlb__sector_hits_T_21;
  wire  tlb_hitsVec_2 = tlb_vm_enabled & tlb__hitsVec_T_17;
  wire  tlb__GEN_13 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_3_valid_1 : tlb_sectored_entries_0_3_valid_0;
  wire  tlb__GEN_14 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_3_valid_2 : tlb__GEN_13;
  wire  tlb__GEN_15 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_3_valid_3 : tlb__GEN_14;
  wire  tlb__hitsVec_T_23 = tlb__GEN_15 & tlb__sector_hits_T_29;
  wire  tlb_hitsVec_3 = tlb_vm_enabled & tlb__hitsVec_T_23;
  wire  tlb__GEN_17 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_4_valid_1 : tlb_sectored_entries_0_4_valid_0;
  wire  tlb__GEN_18 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_4_valid_2 : tlb__GEN_17;
  wire  tlb__GEN_19 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_4_valid_3 : tlb__GEN_18;
  wire  tlb__hitsVec_T_29 = tlb__GEN_19 & tlb__sector_hits_T_37;
  wire  tlb_hitsVec_4 = tlb_vm_enabled & tlb__hitsVec_T_29;
  wire  tlb__GEN_21 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_5_valid_1 : tlb_sectored_entries_0_5_valid_0;
  wire  tlb__GEN_22 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_5_valid_2 : tlb__GEN_21;
  wire  tlb__GEN_23 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_5_valid_3 : tlb__GEN_22;
  wire  tlb__hitsVec_T_35 = tlb__GEN_23 & tlb__sector_hits_T_45;
  wire  tlb_hitsVec_5 = tlb_vm_enabled & tlb__hitsVec_T_35;
  wire  tlb__GEN_25 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_6_valid_1 : tlb_sectored_entries_0_6_valid_0;
  wire  tlb__GEN_26 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_6_valid_2 : tlb__GEN_25;
  wire  tlb__GEN_27 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_6_valid_3 : tlb__GEN_26;
  wire  tlb__hitsVec_T_41 = tlb__GEN_27 & tlb__sector_hits_T_53;
  wire  tlb_hitsVec_6 = tlb_vm_enabled & tlb__hitsVec_T_41;
  wire  tlb__GEN_29 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_7_valid_1 : tlb_sectored_entries_0_7_valid_0;
  wire  tlb__GEN_30 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_7_valid_2 : tlb__GEN_29;
  wire  tlb__GEN_31 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_7_valid_3 : tlb__GEN_30;
  wire  tlb__hitsVec_T_47 = tlb__GEN_31 & tlb__sector_hits_T_61;
  wire  tlb_hitsVec_7 = tlb_vm_enabled & tlb__hitsVec_T_47;
  wire  tlb_hitsVec_8 = tlb_vm_enabled & tlb__superpage_hits_T_4;
  wire  tlb_hitsVec_9 = tlb_vm_enabled & tlb__superpage_hits_T_13;
  wire  tlb_hitsVec_10 = tlb_vm_enabled & tlb__superpage_hits_T_22;
  wire  tlb_hitsVec_11 = tlb_vm_enabled & tlb__superpage_hits_T_31;
  wire [19:0] tlb__hitsVec_T_88 = tlb_special_entry_tag_vpn ^ tlb_vpn;
  wire [9:0] tlb__hitsVec_T_89 = tlb__hitsVec_T_88[19:10];
  wire  tlb__hitsVec_T_90 = tlb__hitsVec_T_89 == 10'h0;
  wire  tlb__hitsVec_T_92 = tlb_special_entry_valid_0 & tlb__hitsVec_T_90;
  wire [9:0] tlb__hitsVec_T_94 = tlb__hitsVec_T_88[9:0];
  wire  tlb__hitsVec_T_95 = tlb__hitsVec_T_94 == 10'h0;
  wire  tlb__hitsVec_T_96 = tlb__mpu_ppn_ignore_T | tlb__hitsVec_T_95;
  wire  tlb__hitsVec_T_97 = tlb__hitsVec_T_92 & tlb__hitsVec_T_96;
  wire  tlb_hitsVec_12 = tlb_vm_enabled & tlb__hitsVec_T_97;
  wire [5:0] tlb_real_hits_lo = {tlb_hitsVec_5,tlb_hitsVec_4,tlb_hitsVec_3,tlb_hitsVec_2,tlb_hitsVec_1,tlb_hitsVec_0};
  wire [12:0] tlb_real_hits = {tlb_hitsVec_12,tlb_hitsVec_11,tlb_hitsVec_10,tlb_hitsVec_9,tlb_hitsVec_8,tlb_hitsVec_7,
    tlb_hitsVec_6,tlb_real_hits_lo};
  wire  tlb__hits_T = ~tlb_vm_enabled;
  wire [13:0] tlb_hits = {tlb__hits_T,tlb_hitsVec_12,tlb_hitsVec_11,tlb_hitsVec_10,tlb_hitsVec_9,tlb_hitsVec_8,
    tlb_hitsVec_7,tlb_hitsVec_6,tlb_real_hits_lo};
  wire  tlb__newEntry_g_T = tlb_io_ptw_resp_bits_pte_g & tlb_io_ptw_resp_bits_pte_v;
  wire  tlb__newEntry_sr_T = ~tlb_io_ptw_resp_bits_pte_w;
  wire  tlb__newEntry_sr_T_1 = tlb_io_ptw_resp_bits_pte_x & tlb__newEntry_sr_T;
  wire  tlb__newEntry_sr_T_2 = tlb_io_ptw_resp_bits_pte_r | tlb__newEntry_sr_T_1;
  wire  tlb__newEntry_sr_T_3 = tlb_io_ptw_resp_bits_pte_v & tlb__newEntry_sr_T_2;
  wire  tlb__newEntry_sr_T_4 = tlb__newEntry_sr_T_3 & tlb_io_ptw_resp_bits_pte_a;
  wire  tlb__newEntry_sr_T_5 = tlb__newEntry_sr_T_4 & tlb_io_ptw_resp_bits_pte_r;
  wire  tlb__newEntry_sw_T_5 = tlb__newEntry_sr_T_4 & tlb_io_ptw_resp_bits_pte_w;
  wire  tlb__newEntry_sw_T_6 = tlb__newEntry_sw_T_5 & tlb_io_ptw_resp_bits_pte_d;
  wire  tlb__newEntry_sx_T_5 = tlb__newEntry_sr_T_4 & tlb_io_ptw_resp_bits_pte_x;
  wire  tlb__T = ~tlb_io_ptw_resp_bits_homogeneous;
  wire [10:0] tlb_special_entry_data_0_lo = {2'h3,tlb_prot_w,tlb_prot_x,tlb_prot_r,tlb__prot_w_T_43,tlb_prot_al,
    tlb_prot_al,tlb_prot_eff,tlb__cacheable_T_49,1'h0};
  wire [4:0] tlb_special_entry_data_0_hi_lo = {1'h0,tlb__newEntry_sw_T_6,tlb__newEntry_sx_T_5,tlb__newEntry_sr_T_5,1'h1}
    ;
  wire [40:0] tlb__special_entry_data_0_T = {tlb_refill_ppn,tlb_io_ptw_resp_bits_pte_u,tlb__newEntry_g_T,
    tlb_io_ptw_resp_bits_ae_ptw,tlb_io_ptw_resp_bits_ae_final,tlb_io_ptw_resp_bits_pf,tlb_special_entry_data_0_hi_lo,
    tlb_special_entry_data_0_lo};
  wire  tlb__T_2 = tlb_io_ptw_resp_bits_level < 1'h1;
  wire  tlb__T_3 = tlb_r_superpage_repl_addr == 2'h0;
  wire  tlb__GEN_32 = tlb_invalidate_refill ? 1'h0 : 1'h1;
  wire  tlb__GEN_36 = tlb__T_3 ? tlb__GEN_32 : tlb_superpage_entries_0_valid_0;
  wire  tlb__T_4 = tlb_r_superpage_repl_addr == 2'h1;
  wire  tlb__GEN_41 = tlb__T_4 ? tlb__GEN_32 : tlb_superpage_entries_1_valid_0;
  wire  tlb__T_5 = tlb_r_superpage_repl_addr == 2'h2;
  wire  tlb__GEN_46 = tlb__T_5 ? tlb__GEN_32 : tlb_superpage_entries_2_valid_0;
  wire  tlb__T_6 = tlb_r_superpage_repl_addr == 2'h3;
  wire  tlb__GEN_51 = tlb__T_6 ? tlb__GEN_32 : tlb_superpage_entries_3_valid_0;
  wire [2:0] tlb_waddr_1 = tlb_r_sectored_hit_valid ? tlb_r_sectored_hit_bits : tlb_r_sectored_repl_addr;
  wire  tlb__T_7 = tlb_waddr_1 == 3'h0;
  wire  tlb__T_8 = ~tlb_r_sectored_hit_valid;
  wire  tlb__GEN_53 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_0_valid_0;
  wire  tlb__GEN_54 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_0_valid_1;
  wire  tlb__GEN_55 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_0_valid_2;
  wire  tlb__GEN_56 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_0_valid_3;
  wire [1:0] tlb_idx = tlb_r_refill_tag[1:0];
  wire  tlb__GEN_57 = 2'h0 == tlb_idx | tlb__GEN_53;
  wire  tlb__GEN_58 = 2'h1 == tlb_idx | tlb__GEN_54;
  wire  tlb__GEN_59 = 2'h2 == tlb_idx | tlb__GEN_55;
  wire  tlb__GEN_60 = 2'h3 == tlb_idx | tlb__GEN_56;
  wire [40:0] tlb__GEN_61 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_0_data_0;
  wire [40:0] tlb__GEN_62 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_0_data_1;
  wire [40:0] tlb__GEN_63 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_0_data_2;
  wire [40:0] tlb__GEN_64 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_0_data_3;
  wire  tlb__GEN_65 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_57;
  wire  tlb__GEN_66 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_58;
  wire  tlb__GEN_67 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_59;
  wire  tlb__GEN_68 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_60;
  wire  tlb__GEN_69 = tlb__T_7 ? tlb__GEN_65 : tlb_sectored_entries_0_0_valid_0;
  wire  tlb__GEN_70 = tlb__T_7 ? tlb__GEN_66 : tlb_sectored_entries_0_0_valid_1;
  wire  tlb__GEN_71 = tlb__T_7 ? tlb__GEN_67 : tlb_sectored_entries_0_0_valid_2;
  wire  tlb__GEN_72 = tlb__T_7 ? tlb__GEN_68 : tlb_sectored_entries_0_0_valid_3;
  wire  tlb__T_9 = tlb_waddr_1 == 3'h1;
  wire  tlb__GEN_80 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_1_valid_0;
  wire  tlb__GEN_81 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_1_valid_1;
  wire  tlb__GEN_82 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_1_valid_2;
  wire  tlb__GEN_83 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_1_valid_3;
  wire  tlb__GEN_84 = 2'h0 == tlb_idx | tlb__GEN_80;
  wire  tlb__GEN_85 = 2'h1 == tlb_idx | tlb__GEN_81;
  wire  tlb__GEN_86 = 2'h2 == tlb_idx | tlb__GEN_82;
  wire  tlb__GEN_87 = 2'h3 == tlb_idx | tlb__GEN_83;
  wire [40:0] tlb__GEN_88 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_1_data_0;
  wire [40:0] tlb__GEN_89 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_1_data_1;
  wire [40:0] tlb__GEN_90 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_1_data_2;
  wire [40:0] tlb__GEN_91 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_1_data_3;
  wire  tlb__GEN_92 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_84;
  wire  tlb__GEN_93 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_85;
  wire  tlb__GEN_94 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_86;
  wire  tlb__GEN_95 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_87;
  wire  tlb__GEN_96 = tlb__T_9 ? tlb__GEN_92 : tlb_sectored_entries_0_1_valid_0;
  wire  tlb__GEN_97 = tlb__T_9 ? tlb__GEN_93 : tlb_sectored_entries_0_1_valid_1;
  wire  tlb__GEN_98 = tlb__T_9 ? tlb__GEN_94 : tlb_sectored_entries_0_1_valid_2;
  wire  tlb__GEN_99 = tlb__T_9 ? tlb__GEN_95 : tlb_sectored_entries_0_1_valid_3;
  wire  tlb__T_11 = tlb_waddr_1 == 3'h2;
  wire  tlb__GEN_107 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_2_valid_0;
  wire  tlb__GEN_108 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_2_valid_1;
  wire  tlb__GEN_109 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_2_valid_2;
  wire  tlb__GEN_110 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_2_valid_3;
  wire  tlb__GEN_111 = 2'h0 == tlb_idx | tlb__GEN_107;
  wire  tlb__GEN_112 = 2'h1 == tlb_idx | tlb__GEN_108;
  wire  tlb__GEN_113 = 2'h2 == tlb_idx | tlb__GEN_109;
  wire  tlb__GEN_114 = 2'h3 == tlb_idx | tlb__GEN_110;
  wire [40:0] tlb__GEN_115 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_2_data_0;
  wire [40:0] tlb__GEN_116 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_2_data_1;
  wire [40:0] tlb__GEN_117 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_2_data_2;
  wire [40:0] tlb__GEN_118 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_2_data_3;
  wire  tlb__GEN_119 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_111;
  wire  tlb__GEN_120 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_112;
  wire  tlb__GEN_121 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_113;
  wire  tlb__GEN_122 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_114;
  wire  tlb__GEN_123 = tlb__T_11 ? tlb__GEN_119 : tlb_sectored_entries_0_2_valid_0;
  wire  tlb__GEN_124 = tlb__T_11 ? tlb__GEN_120 : tlb_sectored_entries_0_2_valid_1;
  wire  tlb__GEN_125 = tlb__T_11 ? tlb__GEN_121 : tlb_sectored_entries_0_2_valid_2;
  wire  tlb__GEN_126 = tlb__T_11 ? tlb__GEN_122 : tlb_sectored_entries_0_2_valid_3;
  wire  tlb__T_13 = tlb_waddr_1 == 3'h3;
  wire  tlb__GEN_134 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_3_valid_0;
  wire  tlb__GEN_135 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_3_valid_1;
  wire  tlb__GEN_136 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_3_valid_2;
  wire  tlb__GEN_137 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_3_valid_3;
  wire  tlb__GEN_138 = 2'h0 == tlb_idx | tlb__GEN_134;
  wire  tlb__GEN_139 = 2'h1 == tlb_idx | tlb__GEN_135;
  wire  tlb__GEN_140 = 2'h2 == tlb_idx | tlb__GEN_136;
  wire  tlb__GEN_141 = 2'h3 == tlb_idx | tlb__GEN_137;
  wire [40:0] tlb__GEN_142 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_3_data_0;
  wire [40:0] tlb__GEN_143 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_3_data_1;
  wire [40:0] tlb__GEN_144 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_3_data_2;
  wire [40:0] tlb__GEN_145 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_3_data_3;
  wire  tlb__GEN_146 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_138;
  wire  tlb__GEN_147 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_139;
  wire  tlb__GEN_148 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_140;
  wire  tlb__GEN_149 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_141;
  wire  tlb__GEN_150 = tlb__T_13 ? tlb__GEN_146 : tlb_sectored_entries_0_3_valid_0;
  wire  tlb__GEN_151 = tlb__T_13 ? tlb__GEN_147 : tlb_sectored_entries_0_3_valid_1;
  wire  tlb__GEN_152 = tlb__T_13 ? tlb__GEN_148 : tlb_sectored_entries_0_3_valid_2;
  wire  tlb__GEN_153 = tlb__T_13 ? tlb__GEN_149 : tlb_sectored_entries_0_3_valid_3;
  wire  tlb__T_15 = tlb_waddr_1 == 3'h4;
  wire  tlb__GEN_161 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_4_valid_0;
  wire  tlb__GEN_162 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_4_valid_1;
  wire  tlb__GEN_163 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_4_valid_2;
  wire  tlb__GEN_164 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_4_valid_3;
  wire  tlb__GEN_165 = 2'h0 == tlb_idx | tlb__GEN_161;
  wire  tlb__GEN_166 = 2'h1 == tlb_idx | tlb__GEN_162;
  wire  tlb__GEN_167 = 2'h2 == tlb_idx | tlb__GEN_163;
  wire  tlb__GEN_168 = 2'h3 == tlb_idx | tlb__GEN_164;
  wire [40:0] tlb__GEN_169 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_4_data_0;
  wire [40:0] tlb__GEN_170 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_4_data_1;
  wire [40:0] tlb__GEN_171 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_4_data_2;
  wire [40:0] tlb__GEN_172 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_4_data_3;
  wire  tlb__GEN_173 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_165;
  wire  tlb__GEN_174 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_166;
  wire  tlb__GEN_175 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_167;
  wire  tlb__GEN_176 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_168;
  wire  tlb__GEN_177 = tlb__T_15 ? tlb__GEN_173 : tlb_sectored_entries_0_4_valid_0;
  wire  tlb__GEN_178 = tlb__T_15 ? tlb__GEN_174 : tlb_sectored_entries_0_4_valid_1;
  wire  tlb__GEN_179 = tlb__T_15 ? tlb__GEN_175 : tlb_sectored_entries_0_4_valid_2;
  wire  tlb__GEN_180 = tlb__T_15 ? tlb__GEN_176 : tlb_sectored_entries_0_4_valid_3;
  wire  tlb__T_17 = tlb_waddr_1 == 3'h5;
  wire  tlb__GEN_188 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_5_valid_0;
  wire  tlb__GEN_189 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_5_valid_1;
  wire  tlb__GEN_190 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_5_valid_2;
  wire  tlb__GEN_191 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_5_valid_3;
  wire  tlb__GEN_192 = 2'h0 == tlb_idx | tlb__GEN_188;
  wire  tlb__GEN_193 = 2'h1 == tlb_idx | tlb__GEN_189;
  wire  tlb__GEN_194 = 2'h2 == tlb_idx | tlb__GEN_190;
  wire  tlb__GEN_195 = 2'h3 == tlb_idx | tlb__GEN_191;
  wire [40:0] tlb__GEN_196 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_5_data_0;
  wire [40:0] tlb__GEN_197 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_5_data_1;
  wire [40:0] tlb__GEN_198 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_5_data_2;
  wire [40:0] tlb__GEN_199 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_5_data_3;
  wire  tlb__GEN_200 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_192;
  wire  tlb__GEN_201 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_193;
  wire  tlb__GEN_202 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_194;
  wire  tlb__GEN_203 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_195;
  wire  tlb__GEN_204 = tlb__T_17 ? tlb__GEN_200 : tlb_sectored_entries_0_5_valid_0;
  wire  tlb__GEN_205 = tlb__T_17 ? tlb__GEN_201 : tlb_sectored_entries_0_5_valid_1;
  wire  tlb__GEN_206 = tlb__T_17 ? tlb__GEN_202 : tlb_sectored_entries_0_5_valid_2;
  wire  tlb__GEN_207 = tlb__T_17 ? tlb__GEN_203 : tlb_sectored_entries_0_5_valid_3;
  wire  tlb__T_19 = tlb_waddr_1 == 3'h6;
  wire  tlb__GEN_215 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_6_valid_0;
  wire  tlb__GEN_216 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_6_valid_1;
  wire  tlb__GEN_217 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_6_valid_2;
  wire  tlb__GEN_218 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_6_valid_3;
  wire  tlb__GEN_219 = 2'h0 == tlb_idx | tlb__GEN_215;
  wire  tlb__GEN_220 = 2'h1 == tlb_idx | tlb__GEN_216;
  wire  tlb__GEN_221 = 2'h2 == tlb_idx | tlb__GEN_217;
  wire  tlb__GEN_222 = 2'h3 == tlb_idx | tlb__GEN_218;
  wire [40:0] tlb__GEN_223 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_6_data_0;
  wire [40:0] tlb__GEN_224 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_6_data_1;
  wire [40:0] tlb__GEN_225 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_6_data_2;
  wire [40:0] tlb__GEN_226 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_6_data_3;
  wire  tlb__GEN_227 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_219;
  wire  tlb__GEN_228 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_220;
  wire  tlb__GEN_229 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_221;
  wire  tlb__GEN_230 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_222;
  wire  tlb__GEN_231 = tlb__T_19 ? tlb__GEN_227 : tlb_sectored_entries_0_6_valid_0;
  wire  tlb__GEN_232 = tlb__T_19 ? tlb__GEN_228 : tlb_sectored_entries_0_6_valid_1;
  wire  tlb__GEN_233 = tlb__T_19 ? tlb__GEN_229 : tlb_sectored_entries_0_6_valid_2;
  wire  tlb__GEN_234 = tlb__T_19 ? tlb__GEN_230 : tlb_sectored_entries_0_6_valid_3;
  wire  tlb__T_21 = tlb_waddr_1 == 3'h7;
  wire  tlb__GEN_242 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_7_valid_0;
  wire  tlb__GEN_243 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_7_valid_1;
  wire  tlb__GEN_244 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_7_valid_2;
  wire  tlb__GEN_245 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_7_valid_3;
  wire  tlb__GEN_246 = 2'h0 == tlb_idx | tlb__GEN_242;
  wire  tlb__GEN_247 = 2'h1 == tlb_idx | tlb__GEN_243;
  wire  tlb__GEN_248 = 2'h2 == tlb_idx | tlb__GEN_244;
  wire  tlb__GEN_249 = 2'h3 == tlb_idx | tlb__GEN_245;
  wire [40:0] tlb__GEN_250 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_7_data_0;
  wire [40:0] tlb__GEN_251 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_7_data_1;
  wire [40:0] tlb__GEN_252 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_7_data_2;
  wire [40:0] tlb__GEN_253 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_7_data_3;
  wire  tlb__GEN_254 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_246;
  wire  tlb__GEN_255 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_247;
  wire  tlb__GEN_256 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_248;
  wire  tlb__GEN_257 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_249;
  wire  tlb__GEN_258 = tlb__T_21 ? tlb__GEN_254 : tlb_sectored_entries_0_7_valid_0;
  wire  tlb__GEN_259 = tlb__T_21 ? tlb__GEN_255 : tlb_sectored_entries_0_7_valid_1;
  wire  tlb__GEN_260 = tlb__T_21 ? tlb__GEN_256 : tlb_sectored_entries_0_7_valid_2;
  wire  tlb__GEN_261 = tlb__T_21 ? tlb__GEN_257 : tlb_sectored_entries_0_7_valid_3;
  wire  tlb__GEN_272 = tlb__T_2 ? tlb__GEN_36 : tlb_superpage_entries_0_valid_0;
  wire  tlb__GEN_277 = tlb__T_2 ? tlb__GEN_41 : tlb_superpage_entries_1_valid_0;
  wire  tlb__GEN_282 = tlb__T_2 ? tlb__GEN_46 : tlb_superpage_entries_2_valid_0;
  wire  tlb__GEN_287 = tlb__T_2 ? tlb__GEN_51 : tlb_superpage_entries_3_valid_0;
  wire  tlb__GEN_289 = tlb__T_2 ? tlb_sectored_entries_0_0_valid_0 : tlb__GEN_69;
  wire  tlb__GEN_290 = tlb__T_2 ? tlb_sectored_entries_0_0_valid_1 : tlb__GEN_70;
  wire  tlb__GEN_291 = tlb__T_2 ? tlb_sectored_entries_0_0_valid_2 : tlb__GEN_71;
  wire  tlb__GEN_292 = tlb__T_2 ? tlb_sectored_entries_0_0_valid_3 : tlb__GEN_72;
  wire  tlb__GEN_300 = tlb__T_2 ? tlb_sectored_entries_0_1_valid_0 : tlb__GEN_96;
  wire  tlb__GEN_301 = tlb__T_2 ? tlb_sectored_entries_0_1_valid_1 : tlb__GEN_97;
  wire  tlb__GEN_302 = tlb__T_2 ? tlb_sectored_entries_0_1_valid_2 : tlb__GEN_98;
  wire  tlb__GEN_303 = tlb__T_2 ? tlb_sectored_entries_0_1_valid_3 : tlb__GEN_99;
  wire  tlb__GEN_311 = tlb__T_2 ? tlb_sectored_entries_0_2_valid_0 : tlb__GEN_123;
  wire  tlb__GEN_312 = tlb__T_2 ? tlb_sectored_entries_0_2_valid_1 : tlb__GEN_124;
  wire  tlb__GEN_313 = tlb__T_2 ? tlb_sectored_entries_0_2_valid_2 : tlb__GEN_125;
  wire  tlb__GEN_314 = tlb__T_2 ? tlb_sectored_entries_0_2_valid_3 : tlb__GEN_126;
  wire  tlb__GEN_322 = tlb__T_2 ? tlb_sectored_entries_0_3_valid_0 : tlb__GEN_150;
  wire  tlb__GEN_323 = tlb__T_2 ? tlb_sectored_entries_0_3_valid_1 : tlb__GEN_151;
  wire  tlb__GEN_324 = tlb__T_2 ? tlb_sectored_entries_0_3_valid_2 : tlb__GEN_152;
  wire  tlb__GEN_325 = tlb__T_2 ? tlb_sectored_entries_0_3_valid_3 : tlb__GEN_153;
  wire  tlb__GEN_333 = tlb__T_2 ? tlb_sectored_entries_0_4_valid_0 : tlb__GEN_177;
  wire  tlb__GEN_334 = tlb__T_2 ? tlb_sectored_entries_0_4_valid_1 : tlb__GEN_178;
  wire  tlb__GEN_335 = tlb__T_2 ? tlb_sectored_entries_0_4_valid_2 : tlb__GEN_179;
  wire  tlb__GEN_336 = tlb__T_2 ? tlb_sectored_entries_0_4_valid_3 : tlb__GEN_180;
  wire  tlb__GEN_344 = tlb__T_2 ? tlb_sectored_entries_0_5_valid_0 : tlb__GEN_204;
  wire  tlb__GEN_345 = tlb__T_2 ? tlb_sectored_entries_0_5_valid_1 : tlb__GEN_205;
  wire  tlb__GEN_346 = tlb__T_2 ? tlb_sectored_entries_0_5_valid_2 : tlb__GEN_206;
  wire  tlb__GEN_347 = tlb__T_2 ? tlb_sectored_entries_0_5_valid_3 : tlb__GEN_207;
  wire  tlb__GEN_355 = tlb__T_2 ? tlb_sectored_entries_0_6_valid_0 : tlb__GEN_231;
  wire  tlb__GEN_356 = tlb__T_2 ? tlb_sectored_entries_0_6_valid_1 : tlb__GEN_232;
  wire  tlb__GEN_357 = tlb__T_2 ? tlb_sectored_entries_0_6_valid_2 : tlb__GEN_233;
  wire  tlb__GEN_358 = tlb__T_2 ? tlb_sectored_entries_0_6_valid_3 : tlb__GEN_234;
  wire  tlb__GEN_366 = tlb__T_2 ? tlb_sectored_entries_0_7_valid_0 : tlb__GEN_258;
  wire  tlb__GEN_367 = tlb__T_2 ? tlb_sectored_entries_0_7_valid_1 : tlb__GEN_259;
  wire  tlb__GEN_368 = tlb__T_2 ? tlb_sectored_entries_0_7_valid_2 : tlb__GEN_260;
  wire  tlb__GEN_369 = tlb__T_2 ? tlb_sectored_entries_0_7_valid_3 : tlb__GEN_261;
  wire  tlb__GEN_380 = tlb__T | tlb_special_entry_valid_0;
  wire  tlb__GEN_385 = tlb__T ? tlb_superpage_entries_0_valid_0 : tlb__GEN_272;
  wire  tlb__GEN_390 = tlb__T ? tlb_superpage_entries_1_valid_0 : tlb__GEN_277;
  wire  tlb__GEN_395 = tlb__T ? tlb_superpage_entries_2_valid_0 : tlb__GEN_282;
  wire  tlb__GEN_400 = tlb__T ? tlb_superpage_entries_3_valid_0 : tlb__GEN_287;
  wire  tlb__GEN_402 = tlb__T ? tlb_sectored_entries_0_0_valid_0 : tlb__GEN_289;
  wire  tlb__GEN_403 = tlb__T ? tlb_sectored_entries_0_0_valid_1 : tlb__GEN_290;
  wire  tlb__GEN_404 = tlb__T ? tlb_sectored_entries_0_0_valid_2 : tlb__GEN_291;
  wire  tlb__GEN_405 = tlb__T ? tlb_sectored_entries_0_0_valid_3 : tlb__GEN_292;
  wire  tlb__GEN_413 = tlb__T ? tlb_sectored_entries_0_1_valid_0 : tlb__GEN_300;
  wire  tlb__GEN_414 = tlb__T ? tlb_sectored_entries_0_1_valid_1 : tlb__GEN_301;
  wire  tlb__GEN_415 = tlb__T ? tlb_sectored_entries_0_1_valid_2 : tlb__GEN_302;
  wire  tlb__GEN_416 = tlb__T ? tlb_sectored_entries_0_1_valid_3 : tlb__GEN_303;
  wire  tlb__GEN_424 = tlb__T ? tlb_sectored_entries_0_2_valid_0 : tlb__GEN_311;
  wire  tlb__GEN_425 = tlb__T ? tlb_sectored_entries_0_2_valid_1 : tlb__GEN_312;
  wire  tlb__GEN_426 = tlb__T ? tlb_sectored_entries_0_2_valid_2 : tlb__GEN_313;
  wire  tlb__GEN_427 = tlb__T ? tlb_sectored_entries_0_2_valid_3 : tlb__GEN_314;
  wire  tlb__GEN_435 = tlb__T ? tlb_sectored_entries_0_3_valid_0 : tlb__GEN_322;
  wire  tlb__GEN_436 = tlb__T ? tlb_sectored_entries_0_3_valid_1 : tlb__GEN_323;
  wire  tlb__GEN_437 = tlb__T ? tlb_sectored_entries_0_3_valid_2 : tlb__GEN_324;
  wire  tlb__GEN_438 = tlb__T ? tlb_sectored_entries_0_3_valid_3 : tlb__GEN_325;
  wire  tlb__GEN_446 = tlb__T ? tlb_sectored_entries_0_4_valid_0 : tlb__GEN_333;
  wire  tlb__GEN_447 = tlb__T ? tlb_sectored_entries_0_4_valid_1 : tlb__GEN_334;
  wire  tlb__GEN_448 = tlb__T ? tlb_sectored_entries_0_4_valid_2 : tlb__GEN_335;
  wire  tlb__GEN_449 = tlb__T ? tlb_sectored_entries_0_4_valid_3 : tlb__GEN_336;
  wire  tlb__GEN_457 = tlb__T ? tlb_sectored_entries_0_5_valid_0 : tlb__GEN_344;
  wire  tlb__GEN_458 = tlb__T ? tlb_sectored_entries_0_5_valid_1 : tlb__GEN_345;
  wire  tlb__GEN_459 = tlb__T ? tlb_sectored_entries_0_5_valid_2 : tlb__GEN_346;
  wire  tlb__GEN_460 = tlb__T ? tlb_sectored_entries_0_5_valid_3 : tlb__GEN_347;
  wire  tlb__GEN_468 = tlb__T ? tlb_sectored_entries_0_6_valid_0 : tlb__GEN_355;
  wire  tlb__GEN_469 = tlb__T ? tlb_sectored_entries_0_6_valid_1 : tlb__GEN_356;
  wire  tlb__GEN_470 = tlb__T ? tlb_sectored_entries_0_6_valid_2 : tlb__GEN_357;
  wire  tlb__GEN_471 = tlb__T ? tlb_sectored_entries_0_6_valid_3 : tlb__GEN_358;
  wire  tlb__GEN_479 = tlb__T ? tlb_sectored_entries_0_7_valid_0 : tlb__GEN_366;
  wire  tlb__GEN_480 = tlb__T ? tlb_sectored_entries_0_7_valid_1 : tlb__GEN_367;
  wire  tlb__GEN_481 = tlb__T ? tlb_sectored_entries_0_7_valid_2 : tlb__GEN_368;
  wire  tlb__GEN_482 = tlb__T ? tlb_sectored_entries_0_7_valid_3 : tlb__GEN_369;
  wire  tlb__GEN_493 = tlb_io_ptw_resp_valid ? tlb__GEN_380 : tlb_special_entry_valid_0;
  wire  tlb__GEN_498 = tlb_io_ptw_resp_valid ? tlb__GEN_385 : tlb_superpage_entries_0_valid_0;
  wire  tlb__GEN_503 = tlb_io_ptw_resp_valid ? tlb__GEN_390 : tlb_superpage_entries_1_valid_0;
  wire  tlb__GEN_508 = tlb_io_ptw_resp_valid ? tlb__GEN_395 : tlb_superpage_entries_2_valid_0;
  wire  tlb__GEN_513 = tlb_io_ptw_resp_valid ? tlb__GEN_400 : tlb_superpage_entries_3_valid_0;
  wire  tlb__GEN_515 = tlb_io_ptw_resp_valid ? tlb__GEN_402 : tlb_sectored_entries_0_0_valid_0;
  wire  tlb__GEN_516 = tlb_io_ptw_resp_valid ? tlb__GEN_403 : tlb_sectored_entries_0_0_valid_1;
  wire  tlb__GEN_517 = tlb_io_ptw_resp_valid ? tlb__GEN_404 : tlb_sectored_entries_0_0_valid_2;
  wire  tlb__GEN_518 = tlb_io_ptw_resp_valid ? tlb__GEN_405 : tlb_sectored_entries_0_0_valid_3;
  wire  tlb__GEN_526 = tlb_io_ptw_resp_valid ? tlb__GEN_413 : tlb_sectored_entries_0_1_valid_0;
  wire  tlb__GEN_527 = tlb_io_ptw_resp_valid ? tlb__GEN_414 : tlb_sectored_entries_0_1_valid_1;
  wire  tlb__GEN_528 = tlb_io_ptw_resp_valid ? tlb__GEN_415 : tlb_sectored_entries_0_1_valid_2;
  wire  tlb__GEN_529 = tlb_io_ptw_resp_valid ? tlb__GEN_416 : tlb_sectored_entries_0_1_valid_3;
  wire  tlb__GEN_537 = tlb_io_ptw_resp_valid ? tlb__GEN_424 : tlb_sectored_entries_0_2_valid_0;
  wire  tlb__GEN_538 = tlb_io_ptw_resp_valid ? tlb__GEN_425 : tlb_sectored_entries_0_2_valid_1;
  wire  tlb__GEN_539 = tlb_io_ptw_resp_valid ? tlb__GEN_426 : tlb_sectored_entries_0_2_valid_2;
  wire  tlb__GEN_540 = tlb_io_ptw_resp_valid ? tlb__GEN_427 : tlb_sectored_entries_0_2_valid_3;
  wire  tlb__GEN_548 = tlb_io_ptw_resp_valid ? tlb__GEN_435 : tlb_sectored_entries_0_3_valid_0;
  wire  tlb__GEN_549 = tlb_io_ptw_resp_valid ? tlb__GEN_436 : tlb_sectored_entries_0_3_valid_1;
  wire  tlb__GEN_550 = tlb_io_ptw_resp_valid ? tlb__GEN_437 : tlb_sectored_entries_0_3_valid_2;
  wire  tlb__GEN_551 = tlb_io_ptw_resp_valid ? tlb__GEN_438 : tlb_sectored_entries_0_3_valid_3;
  wire  tlb__GEN_559 = tlb_io_ptw_resp_valid ? tlb__GEN_446 : tlb_sectored_entries_0_4_valid_0;
  wire  tlb__GEN_560 = tlb_io_ptw_resp_valid ? tlb__GEN_447 : tlb_sectored_entries_0_4_valid_1;
  wire  tlb__GEN_561 = tlb_io_ptw_resp_valid ? tlb__GEN_448 : tlb_sectored_entries_0_4_valid_2;
  wire  tlb__GEN_562 = tlb_io_ptw_resp_valid ? tlb__GEN_449 : tlb_sectored_entries_0_4_valid_3;
  wire  tlb__GEN_570 = tlb_io_ptw_resp_valid ? tlb__GEN_457 : tlb_sectored_entries_0_5_valid_0;
  wire  tlb__GEN_571 = tlb_io_ptw_resp_valid ? tlb__GEN_458 : tlb_sectored_entries_0_5_valid_1;
  wire  tlb__GEN_572 = tlb_io_ptw_resp_valid ? tlb__GEN_459 : tlb_sectored_entries_0_5_valid_2;
  wire  tlb__GEN_573 = tlb_io_ptw_resp_valid ? tlb__GEN_460 : tlb_sectored_entries_0_5_valid_3;
  wire  tlb__GEN_581 = tlb_io_ptw_resp_valid ? tlb__GEN_468 : tlb_sectored_entries_0_6_valid_0;
  wire  tlb__GEN_582 = tlb_io_ptw_resp_valid ? tlb__GEN_469 : tlb_sectored_entries_0_6_valid_1;
  wire  tlb__GEN_583 = tlb_io_ptw_resp_valid ? tlb__GEN_470 : tlb_sectored_entries_0_6_valid_2;
  wire  tlb__GEN_584 = tlb_io_ptw_resp_valid ? tlb__GEN_471 : tlb_sectored_entries_0_6_valid_3;
  wire  tlb__GEN_592 = tlb_io_ptw_resp_valid ? tlb__GEN_479 : tlb_sectored_entries_0_7_valid_0;
  wire  tlb__GEN_593 = tlb_io_ptw_resp_valid ? tlb__GEN_480 : tlb_sectored_entries_0_7_valid_1;
  wire  tlb__GEN_594 = tlb_io_ptw_resp_valid ? tlb__GEN_481 : tlb_sectored_entries_0_7_valid_2;
  wire  tlb__GEN_595 = tlb_io_ptw_resp_valid ? tlb__GEN_482 : tlb_sectored_entries_0_7_valid_3;
  wire [40:0] tlb__GEN_607 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_0_data_1 : tlb_sectored_entries_0_0_data_0
    ;
  wire [40:0] tlb__GEN_608 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_0_data_2 : tlb__GEN_607;
  wire [40:0] tlb__GEN_609 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_0_data_3 : tlb__GEN_608;
  wire [40:0] tlb__GEN_611 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_1_data_1 : tlb_sectored_entries_0_1_data_0
    ;
  wire [40:0] tlb__GEN_612 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_1_data_2 : tlb__GEN_611;
  wire [40:0] tlb__GEN_613 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_1_data_3 : tlb__GEN_612;
  wire [40:0] tlb__GEN_615 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_2_data_1 : tlb_sectored_entries_0_2_data_0
    ;
  wire [40:0] tlb__GEN_616 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_2_data_2 : tlb__GEN_615;
  wire [40:0] tlb__GEN_617 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_2_data_3 : tlb__GEN_616;
  wire [40:0] tlb__GEN_619 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_3_data_1 : tlb_sectored_entries_0_3_data_0
    ;
  wire [40:0] tlb__GEN_620 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_3_data_2 : tlb__GEN_619;
  wire [40:0] tlb__GEN_621 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_3_data_3 : tlb__GEN_620;
  wire [40:0] tlb__GEN_623 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_4_data_1 : tlb_sectored_entries_0_4_data_0
    ;
  wire [40:0] tlb__GEN_624 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_4_data_2 : tlb__GEN_623;
  wire [40:0] tlb__GEN_625 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_4_data_3 : tlb__GEN_624;
  wire [40:0] tlb__GEN_627 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_5_data_1 : tlb_sectored_entries_0_5_data_0
    ;
  wire [40:0] tlb__GEN_628 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_5_data_2 : tlb__GEN_627;
  wire [40:0] tlb__GEN_629 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_5_data_3 : tlb__GEN_628;
  wire [40:0] tlb__GEN_631 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_6_data_1 : tlb_sectored_entries_0_6_data_0
    ;
  wire [40:0] tlb__GEN_632 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_6_data_2 : tlb__GEN_631;
  wire [40:0] tlb__GEN_633 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_6_data_3 : tlb__GEN_632;
  wire [40:0] tlb__GEN_635 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_7_data_1 : tlb_sectored_entries_0_7_data_0
    ;
  wire [40:0] tlb__GEN_636 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_7_data_2 : tlb__GEN_635;
  wire [40:0] tlb__GEN_637 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_7_data_3 : tlb__GEN_636;
  wire  tlb__entries_T_203 = tlb_superpage_entries_0_data_0[19];
  wire  tlb__entries_T_225 = tlb_superpage_entries_1_data_0[19];
  wire  tlb__entries_T_247 = tlb_superpage_entries_2_data_0[19];
  wire  tlb__entries_T_269 = tlb_superpage_entries_3_data_0[19];
  wire [9:0] tlb_ppn_res = tlb_entries_barrier_8_io_y_ppn[19:10];
  wire [19:0] tlb__ppn_T_2 = tlb_vpn | tlb_entries_barrier_8_io_y_ppn;
  wire [9:0] tlb__ppn_T_3 = tlb__ppn_T_2[9:0];
  wire [19:0] tlb__ppn_T_4 = {tlb_ppn_res,tlb__ppn_T_3};
  wire [9:0] tlb_ppn_res_1 = tlb_entries_barrier_9_io_y_ppn[19:10];
  wire [19:0] tlb__ppn_T_6 = tlb_vpn | tlb_entries_barrier_9_io_y_ppn;
  wire [9:0] tlb__ppn_T_7 = tlb__ppn_T_6[9:0];
  wire [19:0] tlb__ppn_T_8 = {tlb_ppn_res_1,tlb__ppn_T_7};
  wire [9:0] tlb_ppn_res_2 = tlb_entries_barrier_10_io_y_ppn[19:10];
  wire [19:0] tlb__ppn_T_10 = tlb_vpn | tlb_entries_barrier_10_io_y_ppn;
  wire [9:0] tlb__ppn_T_11 = tlb__ppn_T_10[9:0];
  wire [19:0] tlb__ppn_T_12 = {tlb_ppn_res_2,tlb__ppn_T_11};
  wire [9:0] tlb_ppn_res_3 = tlb_entries_barrier_11_io_y_ppn[19:10];
  wire [19:0] tlb__ppn_T_14 = tlb_vpn | tlb_entries_barrier_11_io_y_ppn;
  wire [9:0] tlb__ppn_T_15 = tlb__ppn_T_14[9:0];
  wire [19:0] tlb__ppn_T_16 = {tlb_ppn_res_3,tlb__ppn_T_15};
  wire [9:0] tlb_ppn_res_4 = tlb_entries_barrier_12_io_y_ppn[19:10];
  wire [19:0] tlb__ppn_T_18 = tlb__mpu_ppn_T_23 | tlb_entries_barrier_12_io_y_ppn;
  wire [9:0] tlb__ppn_T_19 = tlb__ppn_T_18[9:0];
  wire [19:0] tlb__ppn_T_20 = {tlb_ppn_res_4,tlb__ppn_T_19};
  wire [19:0] tlb__ppn_T_22 = tlb_hitsVec_0 ? tlb_entries_barrier_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_23 = tlb_hitsVec_1 ? tlb_entries_barrier_1_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_24 = tlb_hitsVec_2 ? tlb_entries_barrier_2_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_25 = tlb_hitsVec_3 ? tlb_entries_barrier_3_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_26 = tlb_hitsVec_4 ? tlb_entries_barrier_4_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_27 = tlb_hitsVec_5 ? tlb_entries_barrier_5_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_28 = tlb_hitsVec_6 ? tlb_entries_barrier_6_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_29 = tlb_hitsVec_7 ? tlb_entries_barrier_7_io_y_ppn : 20'h0;
  wire [19:0] tlb__ppn_T_30 = tlb_hitsVec_8 ? tlb__ppn_T_4 : 20'h0;
  wire [19:0] tlb__ppn_T_31 = tlb_hitsVec_9 ? tlb__ppn_T_8 : 20'h0;
  wire [19:0] tlb__ppn_T_32 = tlb_hitsVec_10 ? tlb__ppn_T_12 : 20'h0;
  wire [19:0] tlb__ppn_T_33 = tlb_hitsVec_11 ? tlb__ppn_T_16 : 20'h0;
  wire [19:0] tlb__ppn_T_34 = tlb_hitsVec_12 ? tlb__ppn_T_20 : 20'h0;
  wire [19:0] tlb__ppn_T_35 = tlb__hits_T ? tlb_vpn : 20'h0;
  wire [19:0] tlb__ppn_T_36 = tlb__ppn_T_22 | tlb__ppn_T_23;
  wire [19:0] tlb__ppn_T_37 = tlb__ppn_T_36 | tlb__ppn_T_24;
  wire [19:0] tlb__ppn_T_38 = tlb__ppn_T_37 | tlb__ppn_T_25;
  wire [19:0] tlb__ppn_T_39 = tlb__ppn_T_38 | tlb__ppn_T_26;
  wire [19:0] tlb__ppn_T_40 = tlb__ppn_T_39 | tlb__ppn_T_27;
  wire [19:0] tlb__ppn_T_41 = tlb__ppn_T_40 | tlb__ppn_T_28;
  wire [19:0] tlb__ppn_T_42 = tlb__ppn_T_41 | tlb__ppn_T_29;
  wire [19:0] tlb__ppn_T_43 = tlb__ppn_T_42 | tlb__ppn_T_30;
  wire [19:0] tlb__ppn_T_44 = tlb__ppn_T_43 | tlb__ppn_T_31;
  wire [19:0] tlb__ppn_T_45 = tlb__ppn_T_44 | tlb__ppn_T_32;
  wire [19:0] tlb__ppn_T_46 = tlb__ppn_T_45 | tlb__ppn_T_33;
  wire [19:0] tlb__ppn_T_47 = tlb__ppn_T_46 | tlb__ppn_T_34;
  wire [19:0] tlb__ppn_T_48 = tlb__ppn_T_47 | tlb__ppn_T_35;
  wire [5:0] tlb_ptw_ae_array_lo = {tlb_entries_barrier_5_io_y_ae_ptw,tlb_entries_barrier_4_io_y_ae_ptw,
    tlb_entries_barrier_3_io_y_ae_ptw,tlb_entries_barrier_2_io_y_ae_ptw,tlb_entries_barrier_1_io_y_ae_ptw,
    tlb_entries_barrier_io_y_ae_ptw};
  wire [13:0] tlb_ptw_ae_array = {1'h0,tlb_entries_barrier_12_io_y_ae_ptw,tlb_entries_barrier_11_io_y_ae_ptw,
    tlb_entries_barrier_10_io_y_ae_ptw,tlb_entries_barrier_9_io_y_ae_ptw,tlb_entries_barrier_8_io_y_ae_ptw,
    tlb_entries_barrier_7_io_y_ae_ptw,tlb_entries_barrier_6_io_y_ae_ptw,tlb_ptw_ae_array_lo};
  wire [5:0] tlb_final_ae_array_lo = {tlb_entries_barrier_5_io_y_ae_final,tlb_entries_barrier_4_io_y_ae_final,
    tlb_entries_barrier_3_io_y_ae_final,tlb_entries_barrier_2_io_y_ae_final,tlb_entries_barrier_1_io_y_ae_final,
    tlb_entries_barrier_io_y_ae_final};
  wire [13:0] tlb_final_ae_array = {1'h0,tlb_entries_barrier_12_io_y_ae_final,tlb_entries_barrier_11_io_y_ae_final,
    tlb_entries_barrier_10_io_y_ae_final,tlb_entries_barrier_9_io_y_ae_final,tlb_entries_barrier_8_io_y_ae_final,
    tlb_entries_barrier_7_io_y_ae_final,tlb_entries_barrier_6_io_y_ae_final,tlb_final_ae_array_lo};
  wire [5:0] tlb_ptw_pf_array_lo = {tlb_entries_barrier_5_io_y_pf,tlb_entries_barrier_4_io_y_pf,
    tlb_entries_barrier_3_io_y_pf,tlb_entries_barrier_2_io_y_pf,tlb_entries_barrier_1_io_y_pf,
    tlb_entries_barrier_io_y_pf};
  wire [13:0] tlb_ptw_pf_array = {1'h0,tlb_entries_barrier_12_io_y_pf,tlb_entries_barrier_11_io_y_pf,
    tlb_entries_barrier_10_io_y_pf,tlb_entries_barrier_9_io_y_pf,tlb_entries_barrier_8_io_y_pf,
    tlb_entries_barrier_7_io_y_pf,tlb_entries_barrier_6_io_y_pf,tlb_ptw_pf_array_lo};
  wire [5:0] tlb_ptw_gf_array_lo = {tlb_entries_barrier_5_io_y_gf,tlb_entries_barrier_4_io_y_gf,
    tlb_entries_barrier_3_io_y_gf,tlb_entries_barrier_2_io_y_gf,tlb_entries_barrier_1_io_y_gf,
    tlb_entries_barrier_io_y_gf};
  wire [13:0] tlb_ptw_gf_array = {1'h0,tlb_entries_barrier_12_io_y_gf,tlb_entries_barrier_11_io_y_gf,
    tlb_entries_barrier_10_io_y_gf,tlb_entries_barrier_9_io_y_gf,tlb_entries_barrier_8_io_y_gf,
    tlb_entries_barrier_7_io_y_gf,tlb_entries_barrier_6_io_y_gf,tlb_ptw_gf_array_lo};
  wire  tlb__priv_rw_ok_T = ~tlb_priv_s;
  wire  tlb__priv_rw_ok_T_1 = tlb__priv_rw_ok_T | tlb_io_ptw_status_sum;
  wire [5:0] tlb_priv_rw_ok_lo = {tlb_entries_barrier_5_io_y_u,tlb_entries_barrier_4_io_y_u,tlb_entries_barrier_3_io_y_u
    ,tlb_entries_barrier_2_io_y_u,tlb_entries_barrier_1_io_y_u,tlb_entries_barrier_io_y_u};
  wire [12:0] tlb__priv_rw_ok_T_2 = {tlb_entries_barrier_12_io_y_u,tlb_entries_barrier_11_io_y_u,
    tlb_entries_barrier_10_io_y_u,tlb_entries_barrier_9_io_y_u,tlb_entries_barrier_8_io_y_u,tlb_entries_barrier_7_io_y_u
    ,tlb_entries_barrier_6_io_y_u,tlb_priv_rw_ok_lo};
  wire [12:0] tlb__priv_rw_ok_T_3 = tlb__priv_rw_ok_T_1 ? tlb__priv_rw_ok_T_2 : 13'h0;
  wire [12:0] tlb__priv_rw_ok_T_5 = ~tlb__priv_rw_ok_T_2;
  wire [12:0] tlb__priv_rw_ok_T_6 = tlb_priv_s ? tlb__priv_rw_ok_T_5 : 13'h0;
  wire [12:0] tlb_priv_rw_ok = tlb__priv_rw_ok_T_3 | tlb__priv_rw_ok_T_6;
  wire [5:0] tlb_r_array_lo = {tlb_entries_barrier_5_io_y_sr,tlb_entries_barrier_4_io_y_sr,tlb_entries_barrier_3_io_y_sr
    ,tlb_entries_barrier_2_io_y_sr,tlb_entries_barrier_1_io_y_sr,tlb_entries_barrier_io_y_sr};
  wire [12:0] tlb__r_array_T = {tlb_entries_barrier_12_io_y_sr,tlb_entries_barrier_11_io_y_sr,
    tlb_entries_barrier_10_io_y_sr,tlb_entries_barrier_9_io_y_sr,tlb_entries_barrier_8_io_y_sr,
    tlb_entries_barrier_7_io_y_sr,tlb_entries_barrier_6_io_y_sr,tlb_r_array_lo};
  wire [5:0] tlb_r_array_lo_1 = {tlb_entries_barrier_5_io_y_sx,tlb_entries_barrier_4_io_y_sx,
    tlb_entries_barrier_3_io_y_sx,tlb_entries_barrier_2_io_y_sx,tlb_entries_barrier_1_io_y_sx,
    tlb_entries_barrier_io_y_sx};
  wire [12:0] tlb__r_array_T_1 = {tlb_entries_barrier_12_io_y_sx,tlb_entries_barrier_11_io_y_sx,
    tlb_entries_barrier_10_io_y_sx,tlb_entries_barrier_9_io_y_sx,tlb_entries_barrier_8_io_y_sx,
    tlb_entries_barrier_7_io_y_sx,tlb_entries_barrier_6_io_y_sx,tlb_r_array_lo_1};
  wire [12:0] tlb__r_array_T_2 = tlb_io_ptw_status_mxr ? tlb__r_array_T_1 : 13'h0;
  wire [12:0] tlb__r_array_T_3 = tlb__r_array_T | tlb__r_array_T_2;
  wire [12:0] tlb__r_array_T_4 = tlb_priv_rw_ok & tlb__r_array_T_3;
  wire [13:0] tlb_r_array = {1'h1,tlb__r_array_T_4};
  wire [5:0] tlb_w_array_lo = {tlb_entries_barrier_5_io_y_sw,tlb_entries_barrier_4_io_y_sw,tlb_entries_barrier_3_io_y_sw
    ,tlb_entries_barrier_2_io_y_sw,tlb_entries_barrier_1_io_y_sw,tlb_entries_barrier_io_y_sw};
  wire [12:0] tlb__w_array_T = {tlb_entries_barrier_12_io_y_sw,tlb_entries_barrier_11_io_y_sw,
    tlb_entries_barrier_10_io_y_sw,tlb_entries_barrier_9_io_y_sw,tlb_entries_barrier_8_io_y_sw,
    tlb_entries_barrier_7_io_y_sw,tlb_entries_barrier_6_io_y_sw,tlb_w_array_lo};
  wire [12:0] tlb__w_array_T_1 = tlb_priv_rw_ok & tlb__w_array_T;
  wire [13:0] tlb_w_array = {1'h1,tlb__w_array_T_1};
  wire [1:0] tlb__pr_array_T_1 = tlb_prot_r ? 2'h3 : 2'h0;
  wire [5:0] tlb_pr_array_lo = {tlb_entries_barrier_5_io_y_pr,tlb_entries_barrier_4_io_y_pr,
    tlb_entries_barrier_3_io_y_pr,tlb_entries_barrier_2_io_y_pr,tlb_entries_barrier_1_io_y_pr,
    tlb_entries_barrier_io_y_pr};
  wire [13:0] tlb__pr_array_T_3 = {tlb__pr_array_T_1,tlb_entries_barrier_11_io_y_pr,tlb_entries_barrier_10_io_y_pr,
    tlb_entries_barrier_9_io_y_pr,tlb_entries_barrier_8_io_y_pr,tlb_entries_barrier_7_io_y_pr,
    tlb_entries_barrier_6_io_y_pr,tlb_pr_array_lo};
  wire [13:0] tlb__pr_array_T_4 = tlb_ptw_ae_array | tlb_final_ae_array;
  wire [13:0] tlb__pr_array_T_5 = ~tlb__pr_array_T_4;
  wire [13:0] tlb_pr_array = tlb__pr_array_T_3 & tlb__pr_array_T_5;
  wire [1:0] tlb__pw_array_T_1 = tlb_prot_w ? 2'h3 : 2'h0;
  wire [5:0] tlb_pw_array_lo = {tlb_entries_barrier_5_io_y_pw,tlb_entries_barrier_4_io_y_pw,
    tlb_entries_barrier_3_io_y_pw,tlb_entries_barrier_2_io_y_pw,tlb_entries_barrier_1_io_y_pw,
    tlb_entries_barrier_io_y_pw};
  wire [13:0] tlb__pw_array_T_3 = {tlb__pw_array_T_1,tlb_entries_barrier_11_io_y_pw,tlb_entries_barrier_10_io_y_pw,
    tlb_entries_barrier_9_io_y_pw,tlb_entries_barrier_8_io_y_pw,tlb_entries_barrier_7_io_y_pw,
    tlb_entries_barrier_6_io_y_pw,tlb_pw_array_lo};
  wire [13:0] tlb_pw_array = tlb__pw_array_T_3 & tlb__pr_array_T_5;
  wire [1:0] tlb__eff_array_T_1 = tlb_prot_eff ? 2'h3 : 2'h0;
  wire [5:0] tlb_eff_array_lo = {tlb_entries_barrier_5_io_y_eff,tlb_entries_barrier_4_io_y_eff,
    tlb_entries_barrier_3_io_y_eff,tlb_entries_barrier_2_io_y_eff,tlb_entries_barrier_1_io_y_eff,
    tlb_entries_barrier_io_y_eff};
  wire [13:0] tlb_eff_array = {tlb__eff_array_T_1,tlb_entries_barrier_11_io_y_eff,tlb_entries_barrier_10_io_y_eff,
    tlb_entries_barrier_9_io_y_eff,tlb_entries_barrier_8_io_y_eff,tlb_entries_barrier_7_io_y_eff,
    tlb_entries_barrier_6_io_y_eff,tlb_eff_array_lo};
  wire [1:0] tlb__c_array_T_1 = tlb__cacheable_T_49 ? 2'h3 : 2'h0;
  wire [5:0] tlb_c_array_lo = {tlb_entries_barrier_5_io_y_c,tlb_entries_barrier_4_io_y_c,tlb_entries_barrier_3_io_y_c,
    tlb_entries_barrier_2_io_y_c,tlb_entries_barrier_1_io_y_c,tlb_entries_barrier_io_y_c};
  wire [13:0] tlb_c_array = {tlb__c_array_T_1,tlb_entries_barrier_11_io_y_c,tlb_entries_barrier_10_io_y_c,
    tlb_entries_barrier_9_io_y_c,tlb_entries_barrier_8_io_y_c,tlb_entries_barrier_7_io_y_c,tlb_entries_barrier_6_io_y_c,
    tlb_c_array_lo};
  wire [1:0] tlb__ppp_array_T_1 = tlb__prot_w_T_43 ? 2'h3 : 2'h0;
  wire [5:0] tlb_ppp_array_lo = {tlb_entries_barrier_5_io_y_ppp,tlb_entries_barrier_4_io_y_ppp,
    tlb_entries_barrier_3_io_y_ppp,tlb_entries_barrier_2_io_y_ppp,tlb_entries_barrier_1_io_y_ppp,
    tlb_entries_barrier_io_y_ppp};
  wire [13:0] tlb_ppp_array = {tlb__ppp_array_T_1,tlb_entries_barrier_11_io_y_ppp,tlb_entries_barrier_10_io_y_ppp,
    tlb_entries_barrier_9_io_y_ppp,tlb_entries_barrier_8_io_y_ppp,tlb_entries_barrier_7_io_y_ppp,
    tlb_entries_barrier_6_io_y_ppp,tlb_ppp_array_lo};
  wire [1:0] tlb__paa_array_T_1 = tlb_prot_al ? 2'h3 : 2'h0;
  wire [5:0] tlb_paa_array_lo = {tlb_entries_barrier_5_io_y_paa,tlb_entries_barrier_4_io_y_paa,
    tlb_entries_barrier_3_io_y_paa,tlb_entries_barrier_2_io_y_paa,tlb_entries_barrier_1_io_y_paa,
    tlb_entries_barrier_io_y_paa};
  wire [13:0] tlb_paa_array = {tlb__paa_array_T_1,tlb_entries_barrier_11_io_y_paa,tlb_entries_barrier_10_io_y_paa,
    tlb_entries_barrier_9_io_y_paa,tlb_entries_barrier_8_io_y_paa,tlb_entries_barrier_7_io_y_paa,
    tlb_entries_barrier_6_io_y_paa,tlb_paa_array_lo};
  wire [5:0] tlb_pal_array_lo = {tlb_entries_barrier_5_io_y_pal,tlb_entries_barrier_4_io_y_pal,
    tlb_entries_barrier_3_io_y_pal,tlb_entries_barrier_2_io_y_pal,tlb_entries_barrier_1_io_y_pal,
    tlb_entries_barrier_io_y_pal};
  wire [13:0] tlb_pal_array = {tlb__paa_array_T_1,tlb_entries_barrier_11_io_y_pal,tlb_entries_barrier_10_io_y_pal,
    tlb_entries_barrier_9_io_y_pal,tlb_entries_barrier_8_io_y_pal,tlb_entries_barrier_7_io_y_pal,
    tlb_entries_barrier_6_io_y_pal,tlb_pal_array_lo};
  wire [13:0] tlb_ppp_array_if_cached = tlb_ppp_array | tlb_c_array;
  wire [13:0] tlb_paa_array_if_cached = tlb_paa_array | tlb_c_array;
  wire [13:0] tlb_pal_array_if_cached = tlb_pal_array | tlb_c_array;
  wire [3:0] tlb__misaligned_T = 4'h1 << tlb_io_req_bits_size;
  wire [3:0] tlb__misaligned_T_2 = tlb__misaligned_T - 4'h1;
  wire [31:0] _GEN_446 = {{28'd0}, tlb__misaligned_T_2};
  wire [31:0] tlb__misaligned_T_3 = tlb_io_req_bits_vaddr & _GEN_446;
  wire  tlb_misaligned = |tlb__misaligned_T_3;
  wire  tlb__cmd_lrsc_T = tlb_io_req_bits_cmd == 5'h6;
  wire  tlb__cmd_lrsc_T_1 = tlb_io_req_bits_cmd == 5'h7;
  wire  tlb__cmd_lrsc_T_2 = tlb__cmd_lrsc_T | tlb__cmd_lrsc_T_1;
  wire  tlb__cmd_amo_logical_T = tlb_io_req_bits_cmd == 5'h4;
  wire  tlb__cmd_amo_logical_T_1 = tlb_io_req_bits_cmd == 5'h9;
  wire  tlb__cmd_amo_logical_T_2 = tlb_io_req_bits_cmd == 5'ha;
  wire  tlb__cmd_amo_logical_T_3 = tlb_io_req_bits_cmd == 5'hb;
  wire  tlb__cmd_amo_logical_T_4 = tlb__cmd_amo_logical_T | tlb__cmd_amo_logical_T_1;
  wire  tlb__cmd_amo_logical_T_5 = tlb__cmd_amo_logical_T_4 | tlb__cmd_amo_logical_T_2;
  wire  tlb__cmd_amo_logical_T_6 = tlb__cmd_amo_logical_T_5 | tlb__cmd_amo_logical_T_3;
  wire  tlb__cmd_amo_arithmetic_T = tlb_io_req_bits_cmd == 5'h8;
  wire  tlb__cmd_amo_arithmetic_T_1 = tlb_io_req_bits_cmd == 5'hc;
  wire  tlb__cmd_amo_arithmetic_T_2 = tlb_io_req_bits_cmd == 5'hd;
  wire  tlb__cmd_amo_arithmetic_T_3 = tlb_io_req_bits_cmd == 5'he;
  wire  tlb__cmd_amo_arithmetic_T_4 = tlb_io_req_bits_cmd == 5'hf;
  wire  tlb__cmd_amo_arithmetic_T_5 = tlb__cmd_amo_arithmetic_T | tlb__cmd_amo_arithmetic_T_1;
  wire  tlb__cmd_amo_arithmetic_T_6 = tlb__cmd_amo_arithmetic_T_5 | tlb__cmd_amo_arithmetic_T_2;
  wire  tlb__cmd_amo_arithmetic_T_7 = tlb__cmd_amo_arithmetic_T_6 | tlb__cmd_amo_arithmetic_T_3;
  wire  tlb__cmd_amo_arithmetic_T_8 = tlb__cmd_amo_arithmetic_T_7 | tlb__cmd_amo_arithmetic_T_4;
  wire  tlb_cmd_put_partial = tlb_io_req_bits_cmd == 5'h11;
  wire  tlb__cmd_read_T = tlb_io_req_bits_cmd == 5'h0;
  wire  tlb__cmd_read_T_1 = tlb_io_req_bits_cmd == 5'h10;
  wire  tlb__cmd_read_T_4 = tlb__cmd_read_T | tlb__cmd_read_T_1;
  wire  tlb__cmd_read_T_5 = tlb__cmd_read_T_4 | tlb__cmd_lrsc_T;
  wire  tlb__cmd_read_T_6 = tlb__cmd_read_T_5 | tlb__cmd_lrsc_T_1;
  wire  tlb__cmd_read_T_23 = tlb__cmd_amo_logical_T_6 | tlb__cmd_amo_arithmetic_T_8;
  wire  tlb_cmd_read = tlb__cmd_read_T_6 | tlb__cmd_read_T_23;
  wire  tlb__cmd_write_T = tlb_io_req_bits_cmd == 5'h1;
  wire  tlb__cmd_write_T_2 = tlb__cmd_write_T | tlb_cmd_put_partial;
  wire  tlb__cmd_write_T_4 = tlb__cmd_write_T_2 | tlb__cmd_lrsc_T_1;
  wire  tlb_cmd_write = tlb__cmd_write_T_4 | tlb__cmd_read_T_23;
  wire  tlb__cmd_write_perms_T = tlb_io_req_bits_cmd == 5'h5;
  wire  tlb__cmd_write_perms_T_1 = tlb_io_req_bits_cmd == 5'h17;
  wire  tlb__cmd_write_perms_T_2 = tlb__cmd_write_perms_T | tlb__cmd_write_perms_T_1;
  wire  tlb_cmd_write_perms = tlb_cmd_write | tlb__cmd_write_perms_T_2;
  wire [13:0] tlb__ae_array_T = tlb_misaligned ? tlb_eff_array : 14'h0;
  wire [13:0] tlb__ae_array_T_1 = ~tlb_c_array;
  wire [13:0] tlb__ae_array_T_2 = tlb__cmd_lrsc_T_2 ? tlb__ae_array_T_1 : 14'h0;
  wire [13:0] tlb_ae_array = tlb__ae_array_T | tlb__ae_array_T_2;
  wire [13:0] tlb__ae_ld_array_T = ~tlb_pr_array;
  wire [13:0] tlb__ae_ld_array_T_1 = tlb_ae_array | tlb__ae_ld_array_T;
  wire [13:0] tlb_ae_ld_array = tlb_cmd_read ? tlb__ae_ld_array_T_1 : 14'h0;
  wire [13:0] tlb__ae_st_array_T = ~tlb_pw_array;
  wire [13:0] tlb__ae_st_array_T_1 = tlb_ae_array | tlb__ae_st_array_T;
  wire [13:0] tlb__ae_st_array_T_2 = tlb_cmd_write_perms ? tlb__ae_st_array_T_1 : 14'h0;
  wire [13:0] tlb__ae_st_array_T_3 = ~tlb_ppp_array_if_cached;
  wire [13:0] tlb__ae_st_array_T_4 = tlb_cmd_put_partial ? tlb__ae_st_array_T_3 : 14'h0;
  wire [13:0] tlb__ae_st_array_T_5 = tlb__ae_st_array_T_2 | tlb__ae_st_array_T_4;
  wire [13:0] tlb__ae_st_array_T_6 = ~tlb_pal_array_if_cached;
  wire [13:0] tlb__ae_st_array_T_7 = tlb__cmd_amo_logical_T_6 ? tlb__ae_st_array_T_6 : 14'h0;
  wire [13:0] tlb__ae_st_array_T_8 = tlb__ae_st_array_T_5 | tlb__ae_st_array_T_7;
  wire [13:0] tlb__ae_st_array_T_9 = ~tlb_paa_array_if_cached;
  wire [13:0] tlb__ae_st_array_T_10 = tlb__cmd_amo_arithmetic_T_8 ? tlb__ae_st_array_T_9 : 14'h0;
  wire [13:0] tlb_ae_st_array = tlb__ae_st_array_T_8 | tlb__ae_st_array_T_10;
  wire [13:0] tlb__pf_ld_array_T_1 = ~tlb_r_array;
  wire [13:0] tlb__pf_ld_array_T_2 = ~tlb_ptw_ae_array;
  wire [13:0] tlb__pf_ld_array_T_3 = tlb__pf_ld_array_T_1 & tlb__pf_ld_array_T_2;
  wire [13:0] tlb__pf_ld_array_T_4 = tlb__pf_ld_array_T_3 | tlb_ptw_pf_array;
  wire [13:0] tlb__pf_ld_array_T_5 = ~tlb_ptw_gf_array;
  wire [13:0] tlb__pf_ld_array_T_6 = tlb__pf_ld_array_T_4 & tlb__pf_ld_array_T_5;
  wire [13:0] tlb_pf_ld_array = tlb_cmd_read ? tlb__pf_ld_array_T_6 : 14'h0;
  wire [13:0] tlb__pf_st_array_T = ~tlb_w_array;
  wire [13:0] tlb__pf_st_array_T_2 = tlb__pf_st_array_T & tlb__pf_ld_array_T_2;
  wire [13:0] tlb__pf_st_array_T_3 = tlb__pf_st_array_T_2 | tlb_ptw_pf_array;
  wire [13:0] tlb__pf_st_array_T_5 = tlb__pf_st_array_T_3 & tlb__pf_ld_array_T_5;
  wire [13:0] tlb_pf_st_array = tlb_cmd_write_perms ? tlb__pf_st_array_T_5 : 14'h0;
  wire  tlb_tlb_hit_if_not_gpa_miss = |tlb_real_hits;
  wire  tlb__tlb_miss_T_4 = ~tlb_tlb_hit_if_not_gpa_miss;
  wire  tlb_tlb_miss = tlb_vm_enabled & tlb__tlb_miss_T_4;
  reg [6:0] tlb_state_vec_0;
  reg [2:0] tlb_state_reg_1;
  wire  tlb__T_23 = tlb_io_req_valid & tlb_vm_enabled;
  wire  tlb__T_24 = tlb_sector_hits_0 | tlb_sector_hits_1;
  wire  tlb__T_25 = tlb__T_24 | tlb_sector_hits_2;
  wire  tlb__T_26 = tlb__T_25 | tlb_sector_hits_3;
  wire  tlb__T_27 = tlb__T_26 | tlb_sector_hits_4;
  wire  tlb__T_28 = tlb__T_27 | tlb_sector_hits_5;
  wire  tlb__T_29 = tlb__T_28 | tlb_sector_hits_6;
  wire  tlb__T_30 = tlb__T_29 | tlb_sector_hits_7;
  wire [7:0] tlb__T_31 = {tlb_sector_hits_7,tlb_sector_hits_6,tlb_sector_hits_5,tlb_sector_hits_4,tlb_sector_hits_3,
    tlb_sector_hits_2,tlb_sector_hits_1,tlb_sector_hits_0};
  wire [3:0] tlb_hi_1 = tlb__T_31[7:4];
  wire [3:0] tlb_lo_1 = tlb__T_31[3:0];
  wire  tlb__T_32 = |tlb_hi_1;
  wire [3:0] tlb__T_33 = tlb_hi_1 | tlb_lo_1;
  wire [1:0] tlb_hi_2 = tlb__T_33[3:2];
  wire [1:0] tlb_lo_2 = tlb__T_33[1:0];
  wire  tlb__T_34 = |tlb_hi_2;
  wire [1:0] tlb__T_35 = tlb_hi_2 | tlb_lo_2;
  wire  tlb__T_36 = tlb__T_35[1];
  wire [2:0] tlb__T_38 = {tlb__T_32,tlb__T_34,tlb__T_36};
  wire  tlb__state_vec_0_set_left_older_T = tlb__T_38[2];
  wire  tlb_state_vec_0_set_left_older = ~tlb__state_vec_0_set_left_older_T;
  wire [2:0] tlb_state_vec_0_left_subtree_state = tlb_state_vec_0[5:3];
  wire [2:0] tlb_state_vec_0_right_subtree_state = tlb_state_vec_0[2:0];
  wire [1:0] tlb__state_vec_0_T = tlb__T_38[1:0];
  wire  tlb__state_vec_0_set_left_older_T_1 = tlb__state_vec_0_T[1];
  wire  tlb_state_vec_0_set_left_older_1 = ~tlb__state_vec_0_set_left_older_T_1;
  wire  tlb_state_vec_0_left_subtree_state_1 = tlb_state_vec_0_left_subtree_state[1];
  wire  tlb_state_vec_0_right_subtree_state_1 = tlb_state_vec_0_left_subtree_state[0];
  wire  tlb__state_vec_0_T_1 = tlb__state_vec_0_T[0];
  wire  tlb__state_vec_0_T_3 = ~tlb__state_vec_0_T_1;
  wire  tlb__state_vec_0_T_4 = tlb_state_vec_0_set_left_older_1 ? tlb_state_vec_0_left_subtree_state_1 :
    tlb__state_vec_0_T_3;
  wire  tlb__state_vec_0_T_8 = tlb_state_vec_0_set_left_older_1 ? tlb__state_vec_0_T_3 :
    tlb_state_vec_0_right_subtree_state_1;
  wire [2:0] tlb__state_vec_0_T_9 = {tlb_state_vec_0_set_left_older_1,tlb__state_vec_0_T_4,tlb__state_vec_0_T_8};
  wire [2:0] tlb__state_vec_0_T_10 = tlb_state_vec_0_set_left_older ? tlb_state_vec_0_left_subtree_state :
    tlb__state_vec_0_T_9;
  wire  tlb_state_vec_0_left_subtree_state_2 = tlb_state_vec_0_right_subtree_state[1];
  wire  tlb_state_vec_0_right_subtree_state_2 = tlb_state_vec_0_right_subtree_state[0];
  wire  tlb__state_vec_0_T_15 = tlb_state_vec_0_set_left_older_1 ? tlb_state_vec_0_left_subtree_state_2 :
    tlb__state_vec_0_T_3;
  wire  tlb__state_vec_0_T_19 = tlb_state_vec_0_set_left_older_1 ? tlb__state_vec_0_T_3 :
    tlb_state_vec_0_right_subtree_state_2;
  wire [2:0] tlb__state_vec_0_T_20 = {tlb_state_vec_0_set_left_older_1,tlb__state_vec_0_T_15,tlb__state_vec_0_T_19};
  wire [2:0] tlb__state_vec_0_T_21 = tlb_state_vec_0_set_left_older ? tlb__state_vec_0_T_20 :
    tlb_state_vec_0_right_subtree_state;
  wire [6:0] tlb__state_vec_0_T_22 = {tlb_state_vec_0_set_left_older,tlb__state_vec_0_T_10,tlb__state_vec_0_T_21};
  wire  tlb__T_39 = tlb__superpage_hits_T_4 | tlb__superpage_hits_T_13;
  wire  tlb__T_40 = tlb__T_39 | tlb__superpage_hits_T_22;
  wire  tlb__T_41 = tlb__T_40 | tlb__superpage_hits_T_31;
  wire [3:0] tlb__T_42 = {tlb__superpage_hits_T_31,tlb__superpage_hits_T_22,tlb__superpage_hits_T_13,
    tlb__superpage_hits_T_4};
  wire [1:0] tlb_hi_4 = tlb__T_42[3:2];
  wire [1:0] tlb_lo_4 = tlb__T_42[1:0];
  wire  tlb__T_43 = |tlb_hi_4;
  wire [1:0] tlb__T_44 = tlb_hi_4 | tlb_lo_4;
  wire  tlb__T_45 = tlb__T_44[1];
  wire [1:0] tlb__T_46 = {tlb__T_43,tlb__T_45};
  wire  tlb__state_reg_set_left_older_T = tlb__T_46[1];
  wire  tlb_state_reg_set_left_older = ~tlb__state_reg_set_left_older_T;
  wire  tlb_state_reg_left_subtree_state = tlb_state_reg_1[1];
  wire  tlb_state_reg_right_subtree_state = tlb_state_reg_1[0];
  wire  tlb__state_reg_T = tlb__T_46[0];
  wire  tlb__state_reg_T_2 = ~tlb__state_reg_T;
  wire  tlb__state_reg_T_3 = tlb_state_reg_set_left_older ? tlb_state_reg_left_subtree_state : tlb__state_reg_T_2;
  wire  tlb__state_reg_T_7 = tlb_state_reg_set_left_older ? tlb__state_reg_T_2 : tlb_state_reg_right_subtree_state;
  wire [2:0] tlb__state_reg_T_8 = {tlb_state_reg_set_left_older,tlb__state_reg_T_3,tlb__state_reg_T_7};
  wire [5:0] tlb__multipleHits_T = tlb_real_hits[5:0];
  wire [2:0] tlb__multipleHits_T_1 = tlb__multipleHits_T[2:0];
  wire  tlb__multipleHits_T_2 = tlb__multipleHits_T_1[0];
  wire [1:0] tlb__multipleHits_T_3 = tlb__multipleHits_T_1[2:1];
  wire  tlb__multipleHits_T_4 = tlb__multipleHits_T_3[0];
  wire  tlb__multipleHits_T_5 = tlb__multipleHits_T_3[1];
  wire  tlb_multipleHits_rightOne_1 = tlb__multipleHits_T_4 | tlb__multipleHits_T_5;
  wire  tlb__multipleHits_T_7 = tlb__multipleHits_T_4 & tlb__multipleHits_T_5;
  wire  tlb_multipleHits_leftOne_2 = tlb__multipleHits_T_2 | tlb_multipleHits_rightOne_1;
  wire  tlb__multipleHits_T_9 = tlb__multipleHits_T_2 & tlb_multipleHits_rightOne_1;
  wire  tlb_multipleHits_leftTwo = tlb__multipleHits_T_7 | tlb__multipleHits_T_9;
  wire [2:0] tlb__multipleHits_T_10 = tlb__multipleHits_T[5:3];
  wire  tlb__multipleHits_T_11 = tlb__multipleHits_T_10[0];
  wire [1:0] tlb__multipleHits_T_12 = tlb__multipleHits_T_10[2:1];
  wire  tlb__multipleHits_T_13 = tlb__multipleHits_T_12[0];
  wire  tlb__multipleHits_T_14 = tlb__multipleHits_T_12[1];
  wire  tlb_multipleHits_rightOne_3 = tlb__multipleHits_T_13 | tlb__multipleHits_T_14;
  wire  tlb__multipleHits_T_16 = tlb__multipleHits_T_13 & tlb__multipleHits_T_14;
  wire  tlb_multipleHits_rightOne_4 = tlb__multipleHits_T_11 | tlb_multipleHits_rightOne_3;
  wire  tlb__multipleHits_T_18 = tlb__multipleHits_T_11 & tlb_multipleHits_rightOne_3;
  wire  tlb_multipleHits_rightTwo_2 = tlb__multipleHits_T_16 | tlb__multipleHits_T_18;
  wire  tlb_multipleHits_leftOne_5 = tlb_multipleHits_leftOne_2 | tlb_multipleHits_rightOne_4;
  wire  tlb__multipleHits_T_19 = tlb_multipleHits_leftTwo | tlb_multipleHits_rightTwo_2;
  wire  tlb__multipleHits_T_20 = tlb_multipleHits_leftOne_2 & tlb_multipleHits_rightOne_4;
  wire  tlb_multipleHits_leftTwo_1 = tlb__multipleHits_T_19 | tlb__multipleHits_T_20;
  wire [6:0] tlb__multipleHits_T_21 = tlb_real_hits[12:6];
  wire [2:0] tlb__multipleHits_T_22 = tlb__multipleHits_T_21[2:0];
  wire  tlb__multipleHits_T_23 = tlb__multipleHits_T_22[0];
  wire [1:0] tlb__multipleHits_T_24 = tlb__multipleHits_T_22[2:1];
  wire  tlb__multipleHits_T_25 = tlb__multipleHits_T_24[0];
  wire  tlb__multipleHits_T_26 = tlb__multipleHits_T_24[1];
  wire  tlb_multipleHits_rightOne_6 = tlb__multipleHits_T_25 | tlb__multipleHits_T_26;
  wire  tlb__multipleHits_T_28 = tlb__multipleHits_T_25 & tlb__multipleHits_T_26;
  wire  tlb_multipleHits_leftOne_8 = tlb__multipleHits_T_23 | tlb_multipleHits_rightOne_6;
  wire  tlb__multipleHits_T_30 = tlb__multipleHits_T_23 & tlb_multipleHits_rightOne_6;
  wire  tlb_multipleHits_leftTwo_2 = tlb__multipleHits_T_28 | tlb__multipleHits_T_30;
  wire [3:0] tlb__multipleHits_T_31 = tlb__multipleHits_T_21[6:3];
  wire [1:0] tlb__multipleHits_T_32 = tlb__multipleHits_T_31[1:0];
  wire  tlb__multipleHits_T_33 = tlb__multipleHits_T_32[0];
  wire  tlb__multipleHits_T_34 = tlb__multipleHits_T_32[1];
  wire  tlb_multipleHits_leftOne_10 = tlb__multipleHits_T_33 | tlb__multipleHits_T_34;
  wire  tlb__multipleHits_T_36 = tlb__multipleHits_T_33 & tlb__multipleHits_T_34;
  wire [1:0] tlb__multipleHits_T_37 = tlb__multipleHits_T_31[3:2];
  wire  tlb__multipleHits_T_38 = tlb__multipleHits_T_37[0];
  wire  tlb__multipleHits_T_39 = tlb__multipleHits_T_37[1];
  wire  tlb_multipleHits_rightOne_9 = tlb__multipleHits_T_38 | tlb__multipleHits_T_39;
  wire  tlb__multipleHits_T_41 = tlb__multipleHits_T_38 & tlb__multipleHits_T_39;
  wire  tlb_multipleHits_rightOne_10 = tlb_multipleHits_leftOne_10 | tlb_multipleHits_rightOne_9;
  wire  tlb__multipleHits_T_42 = tlb__multipleHits_T_36 | tlb__multipleHits_T_41;
  wire  tlb__multipleHits_T_43 = tlb_multipleHits_leftOne_10 & tlb_multipleHits_rightOne_9;
  wire  tlb_multipleHits_rightTwo_5 = tlb__multipleHits_T_42 | tlb__multipleHits_T_43;
  wire  tlb_multipleHits_rightOne_11 = tlb_multipleHits_leftOne_8 | tlb_multipleHits_rightOne_10;
  wire  tlb__multipleHits_T_44 = tlb_multipleHits_leftTwo_2 | tlb_multipleHits_rightTwo_5;
  wire  tlb__multipleHits_T_45 = tlb_multipleHits_leftOne_8 & tlb_multipleHits_rightOne_10;
  wire  tlb_multipleHits_rightTwo_6 = tlb__multipleHits_T_44 | tlb__multipleHits_T_45;
  wire  tlb__multipleHits_T_47 = tlb_multipleHits_leftTwo_1 | tlb_multipleHits_rightTwo_6;
  wire  tlb__multipleHits_T_48 = tlb_multipleHits_leftOne_5 & tlb_multipleHits_rightOne_11;
  wire  tlb_multipleHits = tlb__multipleHits_T_47 | tlb__multipleHits_T_48;
  wire [13:0] tlb__io_resp_pf_ld_T_1 = tlb_pf_ld_array & tlb_hits;
  wire [13:0] tlb__io_resp_pf_st_T_1 = tlb_pf_st_array & tlb_hits;
  wire [13:0] tlb__io_resp_ae_ld_T = tlb_ae_ld_array & tlb_hits;
  wire [13:0] tlb__io_resp_ae_st_T = tlb_ae_st_array & tlb_hits;
  wire [13:0] tlb__io_resp_cacheable_T = tlb_c_array & tlb_hits;
  wire  tlb__io_resp_miss_T_1 = tlb_io_ptw_resp_valid | tlb_tlb_miss;
  wire  tlb__T_49 = tlb_io_req_ready & tlb_io_req_valid;
  wire  tlb__T_50 = tlb__T_49 & tlb_tlb_miss;
  wire  tlb_r_superpage_repl_addr_left_subtree_older = tlb_state_reg_1[2];
  wire  tlb__r_superpage_repl_addr_T_2 = tlb_r_superpage_repl_addr_left_subtree_older ? tlb_state_reg_left_subtree_state
     : tlb_state_reg_right_subtree_state;
  wire [1:0] tlb__r_superpage_repl_addr_T_3 = {tlb_r_superpage_repl_addr_left_subtree_older,
    tlb__r_superpage_repl_addr_T_2};
  wire [3:0] tlb_r_superpage_repl_addr_valids = {tlb_superpage_entries_3_valid_0,tlb_superpage_entries_2_valid_0,
    tlb_superpage_entries_1_valid_0,tlb_superpage_entries_0_valid_0};
  wire  tlb__r_superpage_repl_addr_T_4 = &tlb_r_superpage_repl_addr_valids;
  wire [3:0] tlb__r_superpage_repl_addr_T_5 = ~tlb_r_superpage_repl_addr_valids;
  wire  tlb__r_superpage_repl_addr_T_6 = tlb__r_superpage_repl_addr_T_5[0];
  wire  tlb__r_superpage_repl_addr_T_7 = tlb__r_superpage_repl_addr_T_5[1];
  wire  tlb__r_superpage_repl_addr_T_8 = tlb__r_superpage_repl_addr_T_5[2];
  wire [1:0] tlb__r_superpage_repl_addr_T_10 = tlb__r_superpage_repl_addr_T_8 ? 2'h2 : 2'h3;
  wire  tlb_r_sectored_repl_addr_left_subtree_older = tlb_state_vec_0[6];
  wire  tlb_r_sectored_repl_addr_left_subtree_older_1 = tlb_state_vec_0_left_subtree_state[2];
  wire  tlb__r_sectored_repl_addr_T_2 = tlb_r_sectored_repl_addr_left_subtree_older_1 ?
    tlb_state_vec_0_left_subtree_state_1 : tlb_state_vec_0_right_subtree_state_1;
  wire [1:0] tlb__r_sectored_repl_addr_T_3 = {tlb_r_sectored_repl_addr_left_subtree_older_1,
    tlb__r_sectored_repl_addr_T_2};
  wire  tlb_r_sectored_repl_addr_left_subtree_older_2 = tlb_state_vec_0_right_subtree_state[2];
  wire  tlb__r_sectored_repl_addr_T_6 = tlb_r_sectored_repl_addr_left_subtree_older_2 ?
    tlb_state_vec_0_left_subtree_state_2 : tlb_state_vec_0_right_subtree_state_2;
  wire [1:0] tlb__r_sectored_repl_addr_T_7 = {tlb_r_sectored_repl_addr_left_subtree_older_2,
    tlb__r_sectored_repl_addr_T_6};
  wire [1:0] tlb__r_sectored_repl_addr_T_8 = tlb_r_sectored_repl_addr_left_subtree_older ? tlb__r_sectored_repl_addr_T_3
     : tlb__r_sectored_repl_addr_T_7;
  wire [2:0] tlb__r_sectored_repl_addr_T_9 = {tlb_r_sectored_repl_addr_left_subtree_older,tlb__r_sectored_repl_addr_T_8}
    ;
  wire [7:0] tlb_r_sectored_repl_addr_valids = {tlb__sector_hits_T_58,tlb__sector_hits_T_50,tlb__sector_hits_T_42,
    tlb__sector_hits_T_34,tlb__sector_hits_T_26,tlb__sector_hits_T_18,tlb__sector_hits_T_10,tlb__sector_hits_T_2};
  wire  tlb__r_sectored_repl_addr_T_10 = &tlb_r_sectored_repl_addr_valids;
  wire [7:0] tlb__r_sectored_repl_addr_T_11 = ~tlb_r_sectored_repl_addr_valids;
  wire  tlb__r_sectored_repl_addr_T_12 = tlb__r_sectored_repl_addr_T_11[0];
  wire  tlb__r_sectored_repl_addr_T_13 = tlb__r_sectored_repl_addr_T_11[1];
  wire  tlb__r_sectored_repl_addr_T_14 = tlb__r_sectored_repl_addr_T_11[2];
  wire  tlb__r_sectored_repl_addr_T_15 = tlb__r_sectored_repl_addr_T_11[3];
  wire  tlb__r_sectored_repl_addr_T_16 = tlb__r_sectored_repl_addr_T_11[4];
  wire  tlb__r_sectored_repl_addr_T_17 = tlb__r_sectored_repl_addr_T_11[5];
  wire  tlb__r_sectored_repl_addr_T_18 = tlb__r_sectored_repl_addr_T_11[6];
  wire [2:0] tlb__r_sectored_repl_addr_T_20 = tlb__r_sectored_repl_addr_T_18 ? 3'h6 : 3'h7;
  wire [2:0] tlb__r_sectored_repl_addr_T_21 = tlb__r_sectored_repl_addr_T_17 ? 3'h5 : tlb__r_sectored_repl_addr_T_20;
  wire [2:0] tlb__r_sectored_repl_addr_T_22 = tlb__r_sectored_repl_addr_T_16 ? 3'h4 : tlb__r_sectored_repl_addr_T_21;
  wire [2:0] tlb__r_sectored_repl_addr_T_23 = tlb__r_sectored_repl_addr_T_15 ? 3'h3 : tlb__r_sectored_repl_addr_T_22;
  wire [2:0] tlb__r_sectored_repl_addr_T_24 = tlb__r_sectored_repl_addr_T_14 ? 3'h2 : tlb__r_sectored_repl_addr_T_23;
  wire [1:0] tlb__GEN_644 = tlb__T_50 ? 2'h1 : tlb_state;
  wire [1:0] tlb__GEN_655 = tlb_io_sfence_valid ? 2'h0 : tlb__GEN_644;
  wire [1:0] tlb__state_T = tlb_io_sfence_valid ? 2'h3 : 2'h2;
  wire [1:0] tlb__GEN_656 = tlb_io_ptw_req_ready ? tlb__state_T : tlb__GEN_655;
  wire  tlb__T_52 = tlb_state == 2'h2;
  wire  tlb__T_53 = tlb__T_52 & tlb_io_sfence_valid;
  wire  tlb__T_54 = ~tlb_io_sfence_bits_rs1;
  wire [19:0] tlb__T_55 = tlb_io_sfence_bits_addr[31:12];
  wire  tlb__T_56 = tlb__T_55 == tlb_vpn;
  wire  tlb__T_57 = tlb__T_54 | tlb__T_56;
  wire  tlb__T_59 = ~tlb_reset;
  wire  tlb__T_60 = ~tlb__T_57;
  wire  tlb__T_68 = tlb_sectored_entries_0_0_data_0[0];
  wire  tlb__T_87 = tlb_sectored_entries_0_0_data_0[19];
  wire  tlb__T_90 = tlb_sectored_entries_0_0_data_1[0];
  wire  tlb__T_109 = tlb_sectored_entries_0_0_data_1[19];
  wire  tlb__T_112 = tlb_sectored_entries_0_0_data_2[0];
  wire  tlb__T_131 = tlb_sectored_entries_0_0_data_2[19];
  wire  tlb__T_134 = tlb_sectored_entries_0_0_data_3[0];
  wire  tlb__T_153 = tlb_sectored_entries_0_0_data_3[19];
  wire  tlb__T_158 = 2'h0 == tlb_hitsVec_idx;
  wire  tlb__GEN_661 = tlb__T_158 ? 1'h0 : tlb__GEN_515;
  wire  tlb__T_162 = 2'h1 == tlb_hitsVec_idx;
  wire  tlb__GEN_662 = tlb__T_162 ? 1'h0 : tlb__GEN_516;
  wire  tlb__T_166 = 2'h2 == tlb_hitsVec_idx;
  wire  tlb__GEN_663 = tlb__T_166 ? 1'h0 : tlb__GEN_517;
  wire  tlb__T_170 = 2'h3 == tlb_hitsVec_idx;
  wire  tlb__GEN_664 = tlb__T_170 ? 1'h0 : tlb__GEN_518;
  wire  tlb__GEN_665 = tlb__sector_hits_T_5 ? tlb__GEN_661 : tlb__GEN_515;
  wire  tlb__GEN_666 = tlb__sector_hits_T_5 ? tlb__GEN_662 : tlb__GEN_516;
  wire  tlb__GEN_667 = tlb__sector_hits_T_5 ? tlb__GEN_663 : tlb__GEN_517;
  wire  tlb__GEN_668 = tlb__sector_hits_T_5 ? tlb__GEN_664 : tlb__GEN_518;
  wire [9:0] tlb__T_173 = tlb__sector_hits_T_3[19:10];
  wire  tlb__T_174 = tlb__T_173 == 10'h0;
  wire  tlb__GEN_669 = tlb__T_68 ? 1'h0 : tlb__GEN_665;
  wire  tlb__GEN_670 = tlb__T_90 ? 1'h0 : tlb__GEN_666;
  wire  tlb__GEN_671 = tlb__T_112 ? 1'h0 : tlb__GEN_667;
  wire  tlb__GEN_672 = tlb__T_134 ? 1'h0 : tlb__GEN_668;
  wire  tlb__T_362 = ~tlb__T_87;
  wire  tlb__GEN_677 = tlb__T_362 ? 1'h0 : tlb__GEN_515;
  wire  tlb__T_365 = ~tlb__T_109;
  wire  tlb__GEN_678 = tlb__T_365 ? 1'h0 : tlb__GEN_516;
  wire  tlb__T_368 = ~tlb__T_131;
  wire  tlb__GEN_679 = tlb__T_368 ? 1'h0 : tlb__GEN_517;
  wire  tlb__T_371 = ~tlb__T_153;
  wire  tlb__GEN_680 = tlb__T_371 ? 1'h0 : tlb__GEN_518;
  wire  tlb__GEN_685 = tlb_io_sfence_bits_rs2 & tlb__GEN_677;
  wire  tlb__GEN_686 = tlb_io_sfence_bits_rs2 & tlb__GEN_678;
  wire  tlb__GEN_687 = tlb_io_sfence_bits_rs2 & tlb__GEN_679;
  wire  tlb__GEN_688 = tlb_io_sfence_bits_rs2 & tlb__GEN_680;
  wire  tlb__T_473 = tlb_sectored_entries_0_1_data_0[0];
  wire  tlb__T_492 = tlb_sectored_entries_0_1_data_0[19];
  wire  tlb__T_495 = tlb_sectored_entries_0_1_data_1[0];
  wire  tlb__T_514 = tlb_sectored_entries_0_1_data_1[19];
  wire  tlb__T_517 = tlb_sectored_entries_0_1_data_2[0];
  wire  tlb__T_536 = tlb_sectored_entries_0_1_data_2[19];
  wire  tlb__T_539 = tlb_sectored_entries_0_1_data_3[0];
  wire  tlb__T_558 = tlb_sectored_entries_0_1_data_3[19];
  wire  tlb__GEN_693 = tlb__T_158 ? 1'h0 : tlb__GEN_526;
  wire  tlb__GEN_694 = tlb__T_162 ? 1'h0 : tlb__GEN_527;
  wire  tlb__GEN_695 = tlb__T_166 ? 1'h0 : tlb__GEN_528;
  wire  tlb__GEN_696 = tlb__T_170 ? 1'h0 : tlb__GEN_529;
  wire  tlb__GEN_697 = tlb__sector_hits_T_13 ? tlb__GEN_693 : tlb__GEN_526;
  wire  tlb__GEN_698 = tlb__sector_hits_T_13 ? tlb__GEN_694 : tlb__GEN_527;
  wire  tlb__GEN_699 = tlb__sector_hits_T_13 ? tlb__GEN_695 : tlb__GEN_528;
  wire  tlb__GEN_700 = tlb__sector_hits_T_13 ? tlb__GEN_696 : tlb__GEN_529;
  wire [9:0] tlb__T_578 = tlb__sector_hits_T_11[19:10];
  wire  tlb__T_579 = tlb__T_578 == 10'h0;
  wire  tlb__GEN_701 = tlb__T_473 ? 1'h0 : tlb__GEN_697;
  wire  tlb__GEN_702 = tlb__T_495 ? 1'h0 : tlb__GEN_698;
  wire  tlb__GEN_703 = tlb__T_517 ? 1'h0 : tlb__GEN_699;
  wire  tlb__GEN_704 = tlb__T_539 ? 1'h0 : tlb__GEN_700;
  wire  tlb__T_767 = ~tlb__T_492;
  wire  tlb__GEN_709 = tlb__T_767 ? 1'h0 : tlb__GEN_526;
  wire  tlb__T_770 = ~tlb__T_514;
  wire  tlb__GEN_710 = tlb__T_770 ? 1'h0 : tlb__GEN_527;
  wire  tlb__T_773 = ~tlb__T_536;
  wire  tlb__GEN_711 = tlb__T_773 ? 1'h0 : tlb__GEN_528;
  wire  tlb__T_776 = ~tlb__T_558;
  wire  tlb__GEN_712 = tlb__T_776 ? 1'h0 : tlb__GEN_529;
  wire  tlb__GEN_717 = tlb_io_sfence_bits_rs2 & tlb__GEN_709;
  wire  tlb__GEN_718 = tlb_io_sfence_bits_rs2 & tlb__GEN_710;
  wire  tlb__GEN_719 = tlb_io_sfence_bits_rs2 & tlb__GEN_711;
  wire  tlb__GEN_720 = tlb_io_sfence_bits_rs2 & tlb__GEN_712;
  wire  tlb__T_878 = tlb_sectored_entries_0_2_data_0[0];
  wire  tlb__T_897 = tlb_sectored_entries_0_2_data_0[19];
  wire  tlb__T_900 = tlb_sectored_entries_0_2_data_1[0];
  wire  tlb__T_919 = tlb_sectored_entries_0_2_data_1[19];
  wire  tlb__T_922 = tlb_sectored_entries_0_2_data_2[0];
  wire  tlb__T_941 = tlb_sectored_entries_0_2_data_2[19];
  wire  tlb__T_944 = tlb_sectored_entries_0_2_data_3[0];
  wire  tlb__T_963 = tlb_sectored_entries_0_2_data_3[19];
  wire  tlb__GEN_725 = tlb__T_158 ? 1'h0 : tlb__GEN_537;
  wire  tlb__GEN_726 = tlb__T_162 ? 1'h0 : tlb__GEN_538;
  wire  tlb__GEN_727 = tlb__T_166 ? 1'h0 : tlb__GEN_539;
  wire  tlb__GEN_728 = tlb__T_170 ? 1'h0 : tlb__GEN_540;
  wire  tlb__GEN_729 = tlb__sector_hits_T_21 ? tlb__GEN_725 : tlb__GEN_537;
  wire  tlb__GEN_730 = tlb__sector_hits_T_21 ? tlb__GEN_726 : tlb__GEN_538;
  wire  tlb__GEN_731 = tlb__sector_hits_T_21 ? tlb__GEN_727 : tlb__GEN_539;
  wire  tlb__GEN_732 = tlb__sector_hits_T_21 ? tlb__GEN_728 : tlb__GEN_540;
  wire [9:0] tlb__T_983 = tlb__sector_hits_T_19[19:10];
  wire  tlb__T_984 = tlb__T_983 == 10'h0;
  wire  tlb__GEN_733 = tlb__T_878 ? 1'h0 : tlb__GEN_729;
  wire  tlb__GEN_734 = tlb__T_900 ? 1'h0 : tlb__GEN_730;
  wire  tlb__GEN_735 = tlb__T_922 ? 1'h0 : tlb__GEN_731;
  wire  tlb__GEN_736 = tlb__T_944 ? 1'h0 : tlb__GEN_732;
  wire  tlb__T_1172 = ~tlb__T_897;
  wire  tlb__GEN_741 = tlb__T_1172 ? 1'h0 : tlb__GEN_537;
  wire  tlb__T_1175 = ~tlb__T_919;
  wire  tlb__GEN_742 = tlb__T_1175 ? 1'h0 : tlb__GEN_538;
  wire  tlb__T_1178 = ~tlb__T_941;
  wire  tlb__GEN_743 = tlb__T_1178 ? 1'h0 : tlb__GEN_539;
  wire  tlb__T_1181 = ~tlb__T_963;
  wire  tlb__GEN_744 = tlb__T_1181 ? 1'h0 : tlb__GEN_540;
  wire  tlb__GEN_749 = tlb_io_sfence_bits_rs2 & tlb__GEN_741;
  wire  tlb__GEN_750 = tlb_io_sfence_bits_rs2 & tlb__GEN_742;
  wire  tlb__GEN_751 = tlb_io_sfence_bits_rs2 & tlb__GEN_743;
  wire  tlb__GEN_752 = tlb_io_sfence_bits_rs2 & tlb__GEN_744;
  wire  tlb__T_1283 = tlb_sectored_entries_0_3_data_0[0];
  wire  tlb__T_1302 = tlb_sectored_entries_0_3_data_0[19];
  wire  tlb__T_1305 = tlb_sectored_entries_0_3_data_1[0];
  wire  tlb__T_1324 = tlb_sectored_entries_0_3_data_1[19];
  wire  tlb__T_1327 = tlb_sectored_entries_0_3_data_2[0];
  wire  tlb__T_1346 = tlb_sectored_entries_0_3_data_2[19];
  wire  tlb__T_1349 = tlb_sectored_entries_0_3_data_3[0];
  wire  tlb__T_1368 = tlb_sectored_entries_0_3_data_3[19];
  wire  tlb__GEN_757 = tlb__T_158 ? 1'h0 : tlb__GEN_548;
  wire  tlb__GEN_758 = tlb__T_162 ? 1'h0 : tlb__GEN_549;
  wire  tlb__GEN_759 = tlb__T_166 ? 1'h0 : tlb__GEN_550;
  wire  tlb__GEN_760 = tlb__T_170 ? 1'h0 : tlb__GEN_551;
  wire  tlb__GEN_761 = tlb__sector_hits_T_29 ? tlb__GEN_757 : tlb__GEN_548;
  wire  tlb__GEN_762 = tlb__sector_hits_T_29 ? tlb__GEN_758 : tlb__GEN_549;
  wire  tlb__GEN_763 = tlb__sector_hits_T_29 ? tlb__GEN_759 : tlb__GEN_550;
  wire  tlb__GEN_764 = tlb__sector_hits_T_29 ? tlb__GEN_760 : tlb__GEN_551;
  wire [9:0] tlb__T_1388 = tlb__sector_hits_T_27[19:10];
  wire  tlb__T_1389 = tlb__T_1388 == 10'h0;
  wire  tlb__GEN_765 = tlb__T_1283 ? 1'h0 : tlb__GEN_761;
  wire  tlb__GEN_766 = tlb__T_1305 ? 1'h0 : tlb__GEN_762;
  wire  tlb__GEN_767 = tlb__T_1327 ? 1'h0 : tlb__GEN_763;
  wire  tlb__GEN_768 = tlb__T_1349 ? 1'h0 : tlb__GEN_764;
  wire  tlb__T_1577 = ~tlb__T_1302;
  wire  tlb__GEN_773 = tlb__T_1577 ? 1'h0 : tlb__GEN_548;
  wire  tlb__T_1580 = ~tlb__T_1324;
  wire  tlb__GEN_774 = tlb__T_1580 ? 1'h0 : tlb__GEN_549;
  wire  tlb__T_1583 = ~tlb__T_1346;
  wire  tlb__GEN_775 = tlb__T_1583 ? 1'h0 : tlb__GEN_550;
  wire  tlb__T_1586 = ~tlb__T_1368;
  wire  tlb__GEN_776 = tlb__T_1586 ? 1'h0 : tlb__GEN_551;
  wire  tlb__GEN_781 = tlb_io_sfence_bits_rs2 & tlb__GEN_773;
  wire  tlb__GEN_782 = tlb_io_sfence_bits_rs2 & tlb__GEN_774;
  wire  tlb__GEN_783 = tlb_io_sfence_bits_rs2 & tlb__GEN_775;
  wire  tlb__GEN_784 = tlb_io_sfence_bits_rs2 & tlb__GEN_776;
  wire  tlb__T_1688 = tlb_sectored_entries_0_4_data_0[0];
  wire  tlb__T_1707 = tlb_sectored_entries_0_4_data_0[19];
  wire  tlb__T_1710 = tlb_sectored_entries_0_4_data_1[0];
  wire  tlb__T_1729 = tlb_sectored_entries_0_4_data_1[19];
  wire  tlb__T_1732 = tlb_sectored_entries_0_4_data_2[0];
  wire  tlb__T_1751 = tlb_sectored_entries_0_4_data_2[19];
  wire  tlb__T_1754 = tlb_sectored_entries_0_4_data_3[0];
  wire  tlb__T_1773 = tlb_sectored_entries_0_4_data_3[19];
  wire  tlb__GEN_789 = tlb__T_158 ? 1'h0 : tlb__GEN_559;
  wire  tlb__GEN_790 = tlb__T_162 ? 1'h0 : tlb__GEN_560;
  wire  tlb__GEN_791 = tlb__T_166 ? 1'h0 : tlb__GEN_561;
  wire  tlb__GEN_792 = tlb__T_170 ? 1'h0 : tlb__GEN_562;
  wire  tlb__GEN_793 = tlb__sector_hits_T_37 ? tlb__GEN_789 : tlb__GEN_559;
  wire  tlb__GEN_794 = tlb__sector_hits_T_37 ? tlb__GEN_790 : tlb__GEN_560;
  wire  tlb__GEN_795 = tlb__sector_hits_T_37 ? tlb__GEN_791 : tlb__GEN_561;
  wire  tlb__GEN_796 = tlb__sector_hits_T_37 ? tlb__GEN_792 : tlb__GEN_562;
  wire [9:0] tlb__T_1793 = tlb__sector_hits_T_35[19:10];
  wire  tlb__T_1794 = tlb__T_1793 == 10'h0;
  wire  tlb__GEN_797 = tlb__T_1688 ? 1'h0 : tlb__GEN_793;
  wire  tlb__GEN_798 = tlb__T_1710 ? 1'h0 : tlb__GEN_794;
  wire  tlb__GEN_799 = tlb__T_1732 ? 1'h0 : tlb__GEN_795;
  wire  tlb__GEN_800 = tlb__T_1754 ? 1'h0 : tlb__GEN_796;
  wire  tlb__T_1982 = ~tlb__T_1707;
  wire  tlb__GEN_805 = tlb__T_1982 ? 1'h0 : tlb__GEN_559;
  wire  tlb__T_1985 = ~tlb__T_1729;
  wire  tlb__GEN_806 = tlb__T_1985 ? 1'h0 : tlb__GEN_560;
  wire  tlb__T_1988 = ~tlb__T_1751;
  wire  tlb__GEN_807 = tlb__T_1988 ? 1'h0 : tlb__GEN_561;
  wire  tlb__T_1991 = ~tlb__T_1773;
  wire  tlb__GEN_808 = tlb__T_1991 ? 1'h0 : tlb__GEN_562;
  wire  tlb__GEN_813 = tlb_io_sfence_bits_rs2 & tlb__GEN_805;
  wire  tlb__GEN_814 = tlb_io_sfence_bits_rs2 & tlb__GEN_806;
  wire  tlb__GEN_815 = tlb_io_sfence_bits_rs2 & tlb__GEN_807;
  wire  tlb__GEN_816 = tlb_io_sfence_bits_rs2 & tlb__GEN_808;
  wire  tlb__T_2093 = tlb_sectored_entries_0_5_data_0[0];
  wire  tlb__T_2112 = tlb_sectored_entries_0_5_data_0[19];
  wire  tlb__T_2115 = tlb_sectored_entries_0_5_data_1[0];
  wire  tlb__T_2134 = tlb_sectored_entries_0_5_data_1[19];
  wire  tlb__T_2137 = tlb_sectored_entries_0_5_data_2[0];
  wire  tlb__T_2156 = tlb_sectored_entries_0_5_data_2[19];
  wire  tlb__T_2159 = tlb_sectored_entries_0_5_data_3[0];
  wire  tlb__T_2178 = tlb_sectored_entries_0_5_data_3[19];
  wire  tlb__GEN_821 = tlb__T_158 ? 1'h0 : tlb__GEN_570;
  wire  tlb__GEN_822 = tlb__T_162 ? 1'h0 : tlb__GEN_571;
  wire  tlb__GEN_823 = tlb__T_166 ? 1'h0 : tlb__GEN_572;
  wire  tlb__GEN_824 = tlb__T_170 ? 1'h0 : tlb__GEN_573;
  wire  tlb__GEN_825 = tlb__sector_hits_T_45 ? tlb__GEN_821 : tlb__GEN_570;
  wire  tlb__GEN_826 = tlb__sector_hits_T_45 ? tlb__GEN_822 : tlb__GEN_571;
  wire  tlb__GEN_827 = tlb__sector_hits_T_45 ? tlb__GEN_823 : tlb__GEN_572;
  wire  tlb__GEN_828 = tlb__sector_hits_T_45 ? tlb__GEN_824 : tlb__GEN_573;
  wire [9:0] tlb__T_2198 = tlb__sector_hits_T_43[19:10];
  wire  tlb__T_2199 = tlb__T_2198 == 10'h0;
  wire  tlb__GEN_829 = tlb__T_2093 ? 1'h0 : tlb__GEN_825;
  wire  tlb__GEN_830 = tlb__T_2115 ? 1'h0 : tlb__GEN_826;
  wire  tlb__GEN_831 = tlb__T_2137 ? 1'h0 : tlb__GEN_827;
  wire  tlb__GEN_832 = tlb__T_2159 ? 1'h0 : tlb__GEN_828;
  wire  tlb__T_2387 = ~tlb__T_2112;
  wire  tlb__GEN_837 = tlb__T_2387 ? 1'h0 : tlb__GEN_570;
  wire  tlb__T_2390 = ~tlb__T_2134;
  wire  tlb__GEN_838 = tlb__T_2390 ? 1'h0 : tlb__GEN_571;
  wire  tlb__T_2393 = ~tlb__T_2156;
  wire  tlb__GEN_839 = tlb__T_2393 ? 1'h0 : tlb__GEN_572;
  wire  tlb__T_2396 = ~tlb__T_2178;
  wire  tlb__GEN_840 = tlb__T_2396 ? 1'h0 : tlb__GEN_573;
  wire  tlb__GEN_845 = tlb_io_sfence_bits_rs2 & tlb__GEN_837;
  wire  tlb__GEN_846 = tlb_io_sfence_bits_rs2 & tlb__GEN_838;
  wire  tlb__GEN_847 = tlb_io_sfence_bits_rs2 & tlb__GEN_839;
  wire  tlb__GEN_848 = tlb_io_sfence_bits_rs2 & tlb__GEN_840;
  wire  tlb__T_2498 = tlb_sectored_entries_0_6_data_0[0];
  wire  tlb__T_2517 = tlb_sectored_entries_0_6_data_0[19];
  wire  tlb__T_2520 = tlb_sectored_entries_0_6_data_1[0];
  wire  tlb__T_2539 = tlb_sectored_entries_0_6_data_1[19];
  wire  tlb__T_2542 = tlb_sectored_entries_0_6_data_2[0];
  wire  tlb__T_2561 = tlb_sectored_entries_0_6_data_2[19];
  wire  tlb__T_2564 = tlb_sectored_entries_0_6_data_3[0];
  wire  tlb__T_2583 = tlb_sectored_entries_0_6_data_3[19];
  wire  tlb__GEN_853 = tlb__T_158 ? 1'h0 : tlb__GEN_581;
  wire  tlb__GEN_854 = tlb__T_162 ? 1'h0 : tlb__GEN_582;
  wire  tlb__GEN_855 = tlb__T_166 ? 1'h0 : tlb__GEN_583;
  wire  tlb__GEN_856 = tlb__T_170 ? 1'h0 : tlb__GEN_584;
  wire  tlb__GEN_857 = tlb__sector_hits_T_53 ? tlb__GEN_853 : tlb__GEN_581;
  wire  tlb__GEN_858 = tlb__sector_hits_T_53 ? tlb__GEN_854 : tlb__GEN_582;
  wire  tlb__GEN_859 = tlb__sector_hits_T_53 ? tlb__GEN_855 : tlb__GEN_583;
  wire  tlb__GEN_860 = tlb__sector_hits_T_53 ? tlb__GEN_856 : tlb__GEN_584;
  wire [9:0] tlb__T_2603 = tlb__sector_hits_T_51[19:10];
  wire  tlb__T_2604 = tlb__T_2603 == 10'h0;
  wire  tlb__GEN_861 = tlb__T_2498 ? 1'h0 : tlb__GEN_857;
  wire  tlb__GEN_862 = tlb__T_2520 ? 1'h0 : tlb__GEN_858;
  wire  tlb__GEN_863 = tlb__T_2542 ? 1'h0 : tlb__GEN_859;
  wire  tlb__GEN_864 = tlb__T_2564 ? 1'h0 : tlb__GEN_860;
  wire  tlb__T_2792 = ~tlb__T_2517;
  wire  tlb__GEN_869 = tlb__T_2792 ? 1'h0 : tlb__GEN_581;
  wire  tlb__T_2795 = ~tlb__T_2539;
  wire  tlb__GEN_870 = tlb__T_2795 ? 1'h0 : tlb__GEN_582;
  wire  tlb__T_2798 = ~tlb__T_2561;
  wire  tlb__GEN_871 = tlb__T_2798 ? 1'h0 : tlb__GEN_583;
  wire  tlb__T_2801 = ~tlb__T_2583;
  wire  tlb__GEN_872 = tlb__T_2801 ? 1'h0 : tlb__GEN_584;
  wire  tlb__GEN_877 = tlb_io_sfence_bits_rs2 & tlb__GEN_869;
  wire  tlb__GEN_878 = tlb_io_sfence_bits_rs2 & tlb__GEN_870;
  wire  tlb__GEN_879 = tlb_io_sfence_bits_rs2 & tlb__GEN_871;
  wire  tlb__GEN_880 = tlb_io_sfence_bits_rs2 & tlb__GEN_872;
  wire  tlb__T_2903 = tlb_sectored_entries_0_7_data_0[0];
  wire  tlb__T_2922 = tlb_sectored_entries_0_7_data_0[19];
  wire  tlb__T_2925 = tlb_sectored_entries_0_7_data_1[0];
  wire  tlb__T_2944 = tlb_sectored_entries_0_7_data_1[19];
  wire  tlb__T_2947 = tlb_sectored_entries_0_7_data_2[0];
  wire  tlb__T_2966 = tlb_sectored_entries_0_7_data_2[19];
  wire  tlb__T_2969 = tlb_sectored_entries_0_7_data_3[0];
  wire  tlb__T_2988 = tlb_sectored_entries_0_7_data_3[19];
  wire  tlb__GEN_885 = tlb__T_158 ? 1'h0 : tlb__GEN_592;
  wire  tlb__GEN_886 = tlb__T_162 ? 1'h0 : tlb__GEN_593;
  wire  tlb__GEN_887 = tlb__T_166 ? 1'h0 : tlb__GEN_594;
  wire  tlb__GEN_888 = tlb__T_170 ? 1'h0 : tlb__GEN_595;
  wire  tlb__GEN_889 = tlb__sector_hits_T_61 ? tlb__GEN_885 : tlb__GEN_592;
  wire  tlb__GEN_890 = tlb__sector_hits_T_61 ? tlb__GEN_886 : tlb__GEN_593;
  wire  tlb__GEN_891 = tlb__sector_hits_T_61 ? tlb__GEN_887 : tlb__GEN_594;
  wire  tlb__GEN_892 = tlb__sector_hits_T_61 ? tlb__GEN_888 : tlb__GEN_595;
  wire [9:0] tlb__T_3008 = tlb__sector_hits_T_59[19:10];
  wire  tlb__T_3009 = tlb__T_3008 == 10'h0;
  wire  tlb__GEN_893 = tlb__T_2903 ? 1'h0 : tlb__GEN_889;
  wire  tlb__GEN_894 = tlb__T_2925 ? 1'h0 : tlb__GEN_890;
  wire  tlb__GEN_895 = tlb__T_2947 ? 1'h0 : tlb__GEN_891;
  wire  tlb__GEN_896 = tlb__T_2969 ? 1'h0 : tlb__GEN_892;
  wire  tlb__T_3197 = ~tlb__T_2922;
  wire  tlb__GEN_901 = tlb__T_3197 ? 1'h0 : tlb__GEN_592;
  wire  tlb__T_3200 = ~tlb__T_2944;
  wire  tlb__GEN_902 = tlb__T_3200 ? 1'h0 : tlb__GEN_593;
  wire  tlb__T_3203 = ~tlb__T_2966;
  wire  tlb__GEN_903 = tlb__T_3203 ? 1'h0 : tlb__GEN_594;
  wire  tlb__T_3206 = ~tlb__T_2988;
  wire  tlb__GEN_904 = tlb__T_3206 ? 1'h0 : tlb__GEN_595;
  wire  tlb__GEN_909 = tlb_io_sfence_bits_rs2 & tlb__GEN_901;
  wire  tlb__GEN_910 = tlb_io_sfence_bits_rs2 & tlb__GEN_902;
  wire  tlb__GEN_911 = tlb_io_sfence_bits_rs2 & tlb__GEN_903;
  wire  tlb__GEN_912 = tlb_io_sfence_bits_rs2 & tlb__GEN_904;
  wire  tlb__T_3338 = ~tlb__entries_T_203;
  wire  tlb__GEN_918 = tlb__T_3338 ? 1'h0 : tlb__GEN_498;
  wire  tlb__GEN_920 = tlb_io_sfence_bits_rs2 & tlb__GEN_918;
  wire  tlb__T_3401 = ~tlb__entries_T_225;
  wire  tlb__GEN_923 = tlb__T_3401 ? 1'h0 : tlb__GEN_503;
  wire  tlb__GEN_925 = tlb_io_sfence_bits_rs2 & tlb__GEN_923;
  wire  tlb__T_3464 = ~tlb__entries_T_247;
  wire  tlb__GEN_928 = tlb__T_3464 ? 1'h0 : tlb__GEN_508;
  wire  tlb__GEN_930 = tlb_io_sfence_bits_rs2 & tlb__GEN_928;
  wire  tlb__T_3527 = ~tlb__entries_T_269;
  wire  tlb__GEN_933 = tlb__T_3527 ? 1'h0 : tlb__GEN_513;
  wire  tlb__GEN_935 = tlb_io_sfence_bits_rs2 & tlb__GEN_933;
  wire  tlb__T_3590 = ~tlb__mpu_ppn_T_20;
  wire  tlb__GEN_938 = tlb__T_3590 ? 1'h0 : tlb__GEN_493;
  wire  tlb__GEN_940 = tlb_io_sfence_bits_rs2 & tlb__GEN_938;
  wire  tlb__T_4470 = tlb_multipleHits | tlb_reset;
  wire [19:0] pma_checker_mpu_ppn_barrier_io_x_ppn;
  wire  pma_checker_mpu_ppn_barrier_io_x_u;
  wire  pma_checker_mpu_ppn_barrier_io_x_ae_ptw;
  wire  pma_checker_mpu_ppn_barrier_io_x_ae_final;
  wire  pma_checker_mpu_ppn_barrier_io_x_pf;
  wire  pma_checker_mpu_ppn_barrier_io_x_gf;
  wire  pma_checker_mpu_ppn_barrier_io_x_sw;
  wire  pma_checker_mpu_ppn_barrier_io_x_sx;
  wire  pma_checker_mpu_ppn_barrier_io_x_sr;
  wire  pma_checker_mpu_ppn_barrier_io_x_pw;
  wire  pma_checker_mpu_ppn_barrier_io_x_px;
  wire  pma_checker_mpu_ppn_barrier_io_x_pr;
  wire  pma_checker_mpu_ppn_barrier_io_x_ppp;
  wire  pma_checker_mpu_ppn_barrier_io_x_pal;
  wire  pma_checker_mpu_ppn_barrier_io_x_paa;
  wire  pma_checker_mpu_ppn_barrier_io_x_eff;
  wire  pma_checker_mpu_ppn_barrier_io_x_c;
  wire [19:0] pma_checker_mpu_ppn_barrier_io_y_ppn;
  wire  pma_checker_mpu_ppn_barrier_io_y_u;
  wire  pma_checker_mpu_ppn_barrier_io_y_ae_ptw;
  wire  pma_checker_mpu_ppn_barrier_io_y_ae_final;
  wire  pma_checker_mpu_ppn_barrier_io_y_pf;
  wire  pma_checker_mpu_ppn_barrier_io_y_gf;
  wire  pma_checker_mpu_ppn_barrier_io_y_sw;
  wire  pma_checker_mpu_ppn_barrier_io_y_sx;
  wire  pma_checker_mpu_ppn_barrier_io_y_sr;
  wire  pma_checker_mpu_ppn_barrier_io_y_pw;
  wire  pma_checker_mpu_ppn_barrier_io_y_px;
  wire  pma_checker_mpu_ppn_barrier_io_y_pr;
  wire  pma_checker_mpu_ppn_barrier_io_y_ppp;
  wire  pma_checker_mpu_ppn_barrier_io_y_pal;
  wire  pma_checker_mpu_ppn_barrier_io_y_paa;
  wire  pma_checker_mpu_ppn_barrier_io_y_eff;
  wire  pma_checker_mpu_ppn_barrier_io_y_c;
  wire [1:0] pma_checker_pmp_io_prv;
  wire  pma_checker_pmp_io_pmp_0_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_0_cfg_a;
  wire  pma_checker_pmp_io_pmp_0_cfg_x;
  wire  pma_checker_pmp_io_pmp_0_cfg_w;
  wire  pma_checker_pmp_io_pmp_0_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_0_addr;
  wire [31:0] pma_checker_pmp_io_pmp_0_mask;
  wire  pma_checker_pmp_io_pmp_1_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_1_cfg_a;
  wire  pma_checker_pmp_io_pmp_1_cfg_x;
  wire  pma_checker_pmp_io_pmp_1_cfg_w;
  wire  pma_checker_pmp_io_pmp_1_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_1_addr;
  wire [31:0] pma_checker_pmp_io_pmp_1_mask;
  wire  pma_checker_pmp_io_pmp_2_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_2_cfg_a;
  wire  pma_checker_pmp_io_pmp_2_cfg_x;
  wire  pma_checker_pmp_io_pmp_2_cfg_w;
  wire  pma_checker_pmp_io_pmp_2_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_2_addr;
  wire [31:0] pma_checker_pmp_io_pmp_2_mask;
  wire  pma_checker_pmp_io_pmp_3_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_3_cfg_a;
  wire  pma_checker_pmp_io_pmp_3_cfg_x;
  wire  pma_checker_pmp_io_pmp_3_cfg_w;
  wire  pma_checker_pmp_io_pmp_3_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_3_addr;
  wire [31:0] pma_checker_pmp_io_pmp_3_mask;
  wire  pma_checker_pmp_io_pmp_4_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_4_cfg_a;
  wire  pma_checker_pmp_io_pmp_4_cfg_x;
  wire  pma_checker_pmp_io_pmp_4_cfg_w;
  wire  pma_checker_pmp_io_pmp_4_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_4_addr;
  wire [31:0] pma_checker_pmp_io_pmp_4_mask;
  wire  pma_checker_pmp_io_pmp_5_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_5_cfg_a;
  wire  pma_checker_pmp_io_pmp_5_cfg_x;
  wire  pma_checker_pmp_io_pmp_5_cfg_w;
  wire  pma_checker_pmp_io_pmp_5_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_5_addr;
  wire [31:0] pma_checker_pmp_io_pmp_5_mask;
  wire  pma_checker_pmp_io_pmp_6_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_6_cfg_a;
  wire  pma_checker_pmp_io_pmp_6_cfg_x;
  wire  pma_checker_pmp_io_pmp_6_cfg_w;
  wire  pma_checker_pmp_io_pmp_6_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_6_addr;
  wire [31:0] pma_checker_pmp_io_pmp_6_mask;
  wire  pma_checker_pmp_io_pmp_7_cfg_l;
  wire [1:0] pma_checker_pmp_io_pmp_7_cfg_a;
  wire  pma_checker_pmp_io_pmp_7_cfg_x;
  wire  pma_checker_pmp_io_pmp_7_cfg_w;
  wire  pma_checker_pmp_io_pmp_7_cfg_r;
  wire [29:0] pma_checker_pmp_io_pmp_7_addr;
  wire [31:0] pma_checker_pmp_io_pmp_7_mask;
  wire [31:0] pma_checker_pmp_io_addr;
  wire  pma_checker_pmp_io_r;
  wire  pma_checker_pmp_io_w;
  wire  pma_checker_pmp_io_x;
  wire [19:0] pma_checker_entries_barrier_io_x_ppn;
  wire  pma_checker_entries_barrier_io_x_u;
  wire  pma_checker_entries_barrier_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_io_x_ae_final;
  wire  pma_checker_entries_barrier_io_x_pf;
  wire  pma_checker_entries_barrier_io_x_gf;
  wire  pma_checker_entries_barrier_io_x_sw;
  wire  pma_checker_entries_barrier_io_x_sx;
  wire  pma_checker_entries_barrier_io_x_sr;
  wire  pma_checker_entries_barrier_io_x_pw;
  wire  pma_checker_entries_barrier_io_x_px;
  wire  pma_checker_entries_barrier_io_x_pr;
  wire  pma_checker_entries_barrier_io_x_ppp;
  wire  pma_checker_entries_barrier_io_x_pal;
  wire  pma_checker_entries_barrier_io_x_paa;
  wire  pma_checker_entries_barrier_io_x_eff;
  wire  pma_checker_entries_barrier_io_x_c;
  wire [19:0] pma_checker_entries_barrier_io_y_ppn;
  wire  pma_checker_entries_barrier_io_y_u;
  wire  pma_checker_entries_barrier_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_io_y_ae_final;
  wire  pma_checker_entries_barrier_io_y_pf;
  wire  pma_checker_entries_barrier_io_y_gf;
  wire  pma_checker_entries_barrier_io_y_sw;
  wire  pma_checker_entries_barrier_io_y_sx;
  wire  pma_checker_entries_barrier_io_y_sr;
  wire  pma_checker_entries_barrier_io_y_pw;
  wire  pma_checker_entries_barrier_io_y_px;
  wire  pma_checker_entries_barrier_io_y_pr;
  wire  pma_checker_entries_barrier_io_y_ppp;
  wire  pma_checker_entries_barrier_io_y_pal;
  wire  pma_checker_entries_barrier_io_y_paa;
  wire  pma_checker_entries_barrier_io_y_eff;
  wire  pma_checker_entries_barrier_io_y_c;
  wire [19:0] pma_checker_entries_barrier_1_io_x_ppn;
  wire  pma_checker_entries_barrier_1_io_x_u;
  wire  pma_checker_entries_barrier_1_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_1_io_x_ae_final;
  wire  pma_checker_entries_barrier_1_io_x_pf;
  wire  pma_checker_entries_barrier_1_io_x_gf;
  wire  pma_checker_entries_barrier_1_io_x_sw;
  wire  pma_checker_entries_barrier_1_io_x_sx;
  wire  pma_checker_entries_barrier_1_io_x_sr;
  wire  pma_checker_entries_barrier_1_io_x_pw;
  wire  pma_checker_entries_barrier_1_io_x_px;
  wire  pma_checker_entries_barrier_1_io_x_pr;
  wire  pma_checker_entries_barrier_1_io_x_ppp;
  wire  pma_checker_entries_barrier_1_io_x_pal;
  wire  pma_checker_entries_barrier_1_io_x_paa;
  wire  pma_checker_entries_barrier_1_io_x_eff;
  wire  pma_checker_entries_barrier_1_io_x_c;
  wire [19:0] pma_checker_entries_barrier_1_io_y_ppn;
  wire  pma_checker_entries_barrier_1_io_y_u;
  wire  pma_checker_entries_barrier_1_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_1_io_y_ae_final;
  wire  pma_checker_entries_barrier_1_io_y_pf;
  wire  pma_checker_entries_barrier_1_io_y_gf;
  wire  pma_checker_entries_barrier_1_io_y_sw;
  wire  pma_checker_entries_barrier_1_io_y_sx;
  wire  pma_checker_entries_barrier_1_io_y_sr;
  wire  pma_checker_entries_barrier_1_io_y_pw;
  wire  pma_checker_entries_barrier_1_io_y_px;
  wire  pma_checker_entries_barrier_1_io_y_pr;
  wire  pma_checker_entries_barrier_1_io_y_ppp;
  wire  pma_checker_entries_barrier_1_io_y_pal;
  wire  pma_checker_entries_barrier_1_io_y_paa;
  wire  pma_checker_entries_barrier_1_io_y_eff;
  wire  pma_checker_entries_barrier_1_io_y_c;
  wire [19:0] pma_checker_entries_barrier_2_io_x_ppn;
  wire  pma_checker_entries_barrier_2_io_x_u;
  wire  pma_checker_entries_barrier_2_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_2_io_x_ae_final;
  wire  pma_checker_entries_barrier_2_io_x_pf;
  wire  pma_checker_entries_barrier_2_io_x_gf;
  wire  pma_checker_entries_barrier_2_io_x_sw;
  wire  pma_checker_entries_barrier_2_io_x_sx;
  wire  pma_checker_entries_barrier_2_io_x_sr;
  wire  pma_checker_entries_barrier_2_io_x_pw;
  wire  pma_checker_entries_barrier_2_io_x_px;
  wire  pma_checker_entries_barrier_2_io_x_pr;
  wire  pma_checker_entries_barrier_2_io_x_ppp;
  wire  pma_checker_entries_barrier_2_io_x_pal;
  wire  pma_checker_entries_barrier_2_io_x_paa;
  wire  pma_checker_entries_barrier_2_io_x_eff;
  wire  pma_checker_entries_barrier_2_io_x_c;
  wire [19:0] pma_checker_entries_barrier_2_io_y_ppn;
  wire  pma_checker_entries_barrier_2_io_y_u;
  wire  pma_checker_entries_barrier_2_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_2_io_y_ae_final;
  wire  pma_checker_entries_barrier_2_io_y_pf;
  wire  pma_checker_entries_barrier_2_io_y_gf;
  wire  pma_checker_entries_barrier_2_io_y_sw;
  wire  pma_checker_entries_barrier_2_io_y_sx;
  wire  pma_checker_entries_barrier_2_io_y_sr;
  wire  pma_checker_entries_barrier_2_io_y_pw;
  wire  pma_checker_entries_barrier_2_io_y_px;
  wire  pma_checker_entries_barrier_2_io_y_pr;
  wire  pma_checker_entries_barrier_2_io_y_ppp;
  wire  pma_checker_entries_barrier_2_io_y_pal;
  wire  pma_checker_entries_barrier_2_io_y_paa;
  wire  pma_checker_entries_barrier_2_io_y_eff;
  wire  pma_checker_entries_barrier_2_io_y_c;
  wire [19:0] pma_checker_entries_barrier_3_io_x_ppn;
  wire  pma_checker_entries_barrier_3_io_x_u;
  wire  pma_checker_entries_barrier_3_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_3_io_x_ae_final;
  wire  pma_checker_entries_barrier_3_io_x_pf;
  wire  pma_checker_entries_barrier_3_io_x_gf;
  wire  pma_checker_entries_barrier_3_io_x_sw;
  wire  pma_checker_entries_barrier_3_io_x_sx;
  wire  pma_checker_entries_barrier_3_io_x_sr;
  wire  pma_checker_entries_barrier_3_io_x_pw;
  wire  pma_checker_entries_barrier_3_io_x_px;
  wire  pma_checker_entries_barrier_3_io_x_pr;
  wire  pma_checker_entries_barrier_3_io_x_ppp;
  wire  pma_checker_entries_barrier_3_io_x_pal;
  wire  pma_checker_entries_barrier_3_io_x_paa;
  wire  pma_checker_entries_barrier_3_io_x_eff;
  wire  pma_checker_entries_barrier_3_io_x_c;
  wire [19:0] pma_checker_entries_barrier_3_io_y_ppn;
  wire  pma_checker_entries_barrier_3_io_y_u;
  wire  pma_checker_entries_barrier_3_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_3_io_y_ae_final;
  wire  pma_checker_entries_barrier_3_io_y_pf;
  wire  pma_checker_entries_barrier_3_io_y_gf;
  wire  pma_checker_entries_barrier_3_io_y_sw;
  wire  pma_checker_entries_barrier_3_io_y_sx;
  wire  pma_checker_entries_barrier_3_io_y_sr;
  wire  pma_checker_entries_barrier_3_io_y_pw;
  wire  pma_checker_entries_barrier_3_io_y_px;
  wire  pma_checker_entries_barrier_3_io_y_pr;
  wire  pma_checker_entries_barrier_3_io_y_ppp;
  wire  pma_checker_entries_barrier_3_io_y_pal;
  wire  pma_checker_entries_barrier_3_io_y_paa;
  wire  pma_checker_entries_barrier_3_io_y_eff;
  wire  pma_checker_entries_barrier_3_io_y_c;
  wire [19:0] pma_checker_entries_barrier_4_io_x_ppn;
  wire  pma_checker_entries_barrier_4_io_x_u;
  wire  pma_checker_entries_barrier_4_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_4_io_x_ae_final;
  wire  pma_checker_entries_barrier_4_io_x_pf;
  wire  pma_checker_entries_barrier_4_io_x_gf;
  wire  pma_checker_entries_barrier_4_io_x_sw;
  wire  pma_checker_entries_barrier_4_io_x_sx;
  wire  pma_checker_entries_barrier_4_io_x_sr;
  wire  pma_checker_entries_barrier_4_io_x_pw;
  wire  pma_checker_entries_barrier_4_io_x_px;
  wire  pma_checker_entries_barrier_4_io_x_pr;
  wire  pma_checker_entries_barrier_4_io_x_ppp;
  wire  pma_checker_entries_barrier_4_io_x_pal;
  wire  pma_checker_entries_barrier_4_io_x_paa;
  wire  pma_checker_entries_barrier_4_io_x_eff;
  wire  pma_checker_entries_barrier_4_io_x_c;
  wire [19:0] pma_checker_entries_barrier_4_io_y_ppn;
  wire  pma_checker_entries_barrier_4_io_y_u;
  wire  pma_checker_entries_barrier_4_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_4_io_y_ae_final;
  wire  pma_checker_entries_barrier_4_io_y_pf;
  wire  pma_checker_entries_barrier_4_io_y_gf;
  wire  pma_checker_entries_barrier_4_io_y_sw;
  wire  pma_checker_entries_barrier_4_io_y_sx;
  wire  pma_checker_entries_barrier_4_io_y_sr;
  wire  pma_checker_entries_barrier_4_io_y_pw;
  wire  pma_checker_entries_barrier_4_io_y_px;
  wire  pma_checker_entries_barrier_4_io_y_pr;
  wire  pma_checker_entries_barrier_4_io_y_ppp;
  wire  pma_checker_entries_barrier_4_io_y_pal;
  wire  pma_checker_entries_barrier_4_io_y_paa;
  wire  pma_checker_entries_barrier_4_io_y_eff;
  wire  pma_checker_entries_barrier_4_io_y_c;
  wire [19:0] pma_checker_entries_barrier_5_io_x_ppn;
  wire  pma_checker_entries_barrier_5_io_x_u;
  wire  pma_checker_entries_barrier_5_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_5_io_x_ae_final;
  wire  pma_checker_entries_barrier_5_io_x_pf;
  wire  pma_checker_entries_barrier_5_io_x_gf;
  wire  pma_checker_entries_barrier_5_io_x_sw;
  wire  pma_checker_entries_barrier_5_io_x_sx;
  wire  pma_checker_entries_barrier_5_io_x_sr;
  wire  pma_checker_entries_barrier_5_io_x_pw;
  wire  pma_checker_entries_barrier_5_io_x_px;
  wire  pma_checker_entries_barrier_5_io_x_pr;
  wire  pma_checker_entries_barrier_5_io_x_ppp;
  wire  pma_checker_entries_barrier_5_io_x_pal;
  wire  pma_checker_entries_barrier_5_io_x_paa;
  wire  pma_checker_entries_barrier_5_io_x_eff;
  wire  pma_checker_entries_barrier_5_io_x_c;
  wire [19:0] pma_checker_entries_barrier_5_io_y_ppn;
  wire  pma_checker_entries_barrier_5_io_y_u;
  wire  pma_checker_entries_barrier_5_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_5_io_y_ae_final;
  wire  pma_checker_entries_barrier_5_io_y_pf;
  wire  pma_checker_entries_barrier_5_io_y_gf;
  wire  pma_checker_entries_barrier_5_io_y_sw;
  wire  pma_checker_entries_barrier_5_io_y_sx;
  wire  pma_checker_entries_barrier_5_io_y_sr;
  wire  pma_checker_entries_barrier_5_io_y_pw;
  wire  pma_checker_entries_barrier_5_io_y_px;
  wire  pma_checker_entries_barrier_5_io_y_pr;
  wire  pma_checker_entries_barrier_5_io_y_ppp;
  wire  pma_checker_entries_barrier_5_io_y_pal;
  wire  pma_checker_entries_barrier_5_io_y_paa;
  wire  pma_checker_entries_barrier_5_io_y_eff;
  wire  pma_checker_entries_barrier_5_io_y_c;
  wire [19:0] pma_checker_entries_barrier_6_io_x_ppn;
  wire  pma_checker_entries_barrier_6_io_x_u;
  wire  pma_checker_entries_barrier_6_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_6_io_x_ae_final;
  wire  pma_checker_entries_barrier_6_io_x_pf;
  wire  pma_checker_entries_barrier_6_io_x_gf;
  wire  pma_checker_entries_barrier_6_io_x_sw;
  wire  pma_checker_entries_barrier_6_io_x_sx;
  wire  pma_checker_entries_barrier_6_io_x_sr;
  wire  pma_checker_entries_barrier_6_io_x_pw;
  wire  pma_checker_entries_barrier_6_io_x_px;
  wire  pma_checker_entries_barrier_6_io_x_pr;
  wire  pma_checker_entries_barrier_6_io_x_ppp;
  wire  pma_checker_entries_barrier_6_io_x_pal;
  wire  pma_checker_entries_barrier_6_io_x_paa;
  wire  pma_checker_entries_barrier_6_io_x_eff;
  wire  pma_checker_entries_barrier_6_io_x_c;
  wire [19:0] pma_checker_entries_barrier_6_io_y_ppn;
  wire  pma_checker_entries_barrier_6_io_y_u;
  wire  pma_checker_entries_barrier_6_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_6_io_y_ae_final;
  wire  pma_checker_entries_barrier_6_io_y_pf;
  wire  pma_checker_entries_barrier_6_io_y_gf;
  wire  pma_checker_entries_barrier_6_io_y_sw;
  wire  pma_checker_entries_barrier_6_io_y_sx;
  wire  pma_checker_entries_barrier_6_io_y_sr;
  wire  pma_checker_entries_barrier_6_io_y_pw;
  wire  pma_checker_entries_barrier_6_io_y_px;
  wire  pma_checker_entries_barrier_6_io_y_pr;
  wire  pma_checker_entries_barrier_6_io_y_ppp;
  wire  pma_checker_entries_barrier_6_io_y_pal;
  wire  pma_checker_entries_barrier_6_io_y_paa;
  wire  pma_checker_entries_barrier_6_io_y_eff;
  wire  pma_checker_entries_barrier_6_io_y_c;
  wire [19:0] pma_checker_entries_barrier_7_io_x_ppn;
  wire  pma_checker_entries_barrier_7_io_x_u;
  wire  pma_checker_entries_barrier_7_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_7_io_x_ae_final;
  wire  pma_checker_entries_barrier_7_io_x_pf;
  wire  pma_checker_entries_barrier_7_io_x_gf;
  wire  pma_checker_entries_barrier_7_io_x_sw;
  wire  pma_checker_entries_barrier_7_io_x_sx;
  wire  pma_checker_entries_barrier_7_io_x_sr;
  wire  pma_checker_entries_barrier_7_io_x_pw;
  wire  pma_checker_entries_barrier_7_io_x_px;
  wire  pma_checker_entries_barrier_7_io_x_pr;
  wire  pma_checker_entries_barrier_7_io_x_ppp;
  wire  pma_checker_entries_barrier_7_io_x_pal;
  wire  pma_checker_entries_barrier_7_io_x_paa;
  wire  pma_checker_entries_barrier_7_io_x_eff;
  wire  pma_checker_entries_barrier_7_io_x_c;
  wire [19:0] pma_checker_entries_barrier_7_io_y_ppn;
  wire  pma_checker_entries_barrier_7_io_y_u;
  wire  pma_checker_entries_barrier_7_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_7_io_y_ae_final;
  wire  pma_checker_entries_barrier_7_io_y_pf;
  wire  pma_checker_entries_barrier_7_io_y_gf;
  wire  pma_checker_entries_barrier_7_io_y_sw;
  wire  pma_checker_entries_barrier_7_io_y_sx;
  wire  pma_checker_entries_barrier_7_io_y_sr;
  wire  pma_checker_entries_barrier_7_io_y_pw;
  wire  pma_checker_entries_barrier_7_io_y_px;
  wire  pma_checker_entries_barrier_7_io_y_pr;
  wire  pma_checker_entries_barrier_7_io_y_ppp;
  wire  pma_checker_entries_barrier_7_io_y_pal;
  wire  pma_checker_entries_barrier_7_io_y_paa;
  wire  pma_checker_entries_barrier_7_io_y_eff;
  wire  pma_checker_entries_barrier_7_io_y_c;
  wire [19:0] pma_checker_entries_barrier_8_io_x_ppn;
  wire  pma_checker_entries_barrier_8_io_x_u;
  wire  pma_checker_entries_barrier_8_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_8_io_x_ae_final;
  wire  pma_checker_entries_barrier_8_io_x_pf;
  wire  pma_checker_entries_barrier_8_io_x_gf;
  wire  pma_checker_entries_barrier_8_io_x_sw;
  wire  pma_checker_entries_barrier_8_io_x_sx;
  wire  pma_checker_entries_barrier_8_io_x_sr;
  wire  pma_checker_entries_barrier_8_io_x_pw;
  wire  pma_checker_entries_barrier_8_io_x_px;
  wire  pma_checker_entries_barrier_8_io_x_pr;
  wire  pma_checker_entries_barrier_8_io_x_ppp;
  wire  pma_checker_entries_barrier_8_io_x_pal;
  wire  pma_checker_entries_barrier_8_io_x_paa;
  wire  pma_checker_entries_barrier_8_io_x_eff;
  wire  pma_checker_entries_barrier_8_io_x_c;
  wire [19:0] pma_checker_entries_barrier_8_io_y_ppn;
  wire  pma_checker_entries_barrier_8_io_y_u;
  wire  pma_checker_entries_barrier_8_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_8_io_y_ae_final;
  wire  pma_checker_entries_barrier_8_io_y_pf;
  wire  pma_checker_entries_barrier_8_io_y_gf;
  wire  pma_checker_entries_barrier_8_io_y_sw;
  wire  pma_checker_entries_barrier_8_io_y_sx;
  wire  pma_checker_entries_barrier_8_io_y_sr;
  wire  pma_checker_entries_barrier_8_io_y_pw;
  wire  pma_checker_entries_barrier_8_io_y_px;
  wire  pma_checker_entries_barrier_8_io_y_pr;
  wire  pma_checker_entries_barrier_8_io_y_ppp;
  wire  pma_checker_entries_barrier_8_io_y_pal;
  wire  pma_checker_entries_barrier_8_io_y_paa;
  wire  pma_checker_entries_barrier_8_io_y_eff;
  wire  pma_checker_entries_barrier_8_io_y_c;
  wire [19:0] pma_checker_entries_barrier_9_io_x_ppn;
  wire  pma_checker_entries_barrier_9_io_x_u;
  wire  pma_checker_entries_barrier_9_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_9_io_x_ae_final;
  wire  pma_checker_entries_barrier_9_io_x_pf;
  wire  pma_checker_entries_barrier_9_io_x_gf;
  wire  pma_checker_entries_barrier_9_io_x_sw;
  wire  pma_checker_entries_barrier_9_io_x_sx;
  wire  pma_checker_entries_barrier_9_io_x_sr;
  wire  pma_checker_entries_barrier_9_io_x_pw;
  wire  pma_checker_entries_barrier_9_io_x_px;
  wire  pma_checker_entries_barrier_9_io_x_pr;
  wire  pma_checker_entries_barrier_9_io_x_ppp;
  wire  pma_checker_entries_barrier_9_io_x_pal;
  wire  pma_checker_entries_barrier_9_io_x_paa;
  wire  pma_checker_entries_barrier_9_io_x_eff;
  wire  pma_checker_entries_barrier_9_io_x_c;
  wire [19:0] pma_checker_entries_barrier_9_io_y_ppn;
  wire  pma_checker_entries_barrier_9_io_y_u;
  wire  pma_checker_entries_barrier_9_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_9_io_y_ae_final;
  wire  pma_checker_entries_barrier_9_io_y_pf;
  wire  pma_checker_entries_barrier_9_io_y_gf;
  wire  pma_checker_entries_barrier_9_io_y_sw;
  wire  pma_checker_entries_barrier_9_io_y_sx;
  wire  pma_checker_entries_barrier_9_io_y_sr;
  wire  pma_checker_entries_barrier_9_io_y_pw;
  wire  pma_checker_entries_barrier_9_io_y_px;
  wire  pma_checker_entries_barrier_9_io_y_pr;
  wire  pma_checker_entries_barrier_9_io_y_ppp;
  wire  pma_checker_entries_barrier_9_io_y_pal;
  wire  pma_checker_entries_barrier_9_io_y_paa;
  wire  pma_checker_entries_barrier_9_io_y_eff;
  wire  pma_checker_entries_barrier_9_io_y_c;
  wire [19:0] pma_checker_entries_barrier_10_io_x_ppn;
  wire  pma_checker_entries_barrier_10_io_x_u;
  wire  pma_checker_entries_barrier_10_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_10_io_x_ae_final;
  wire  pma_checker_entries_barrier_10_io_x_pf;
  wire  pma_checker_entries_barrier_10_io_x_gf;
  wire  pma_checker_entries_barrier_10_io_x_sw;
  wire  pma_checker_entries_barrier_10_io_x_sx;
  wire  pma_checker_entries_barrier_10_io_x_sr;
  wire  pma_checker_entries_barrier_10_io_x_pw;
  wire  pma_checker_entries_barrier_10_io_x_px;
  wire  pma_checker_entries_barrier_10_io_x_pr;
  wire  pma_checker_entries_barrier_10_io_x_ppp;
  wire  pma_checker_entries_barrier_10_io_x_pal;
  wire  pma_checker_entries_barrier_10_io_x_paa;
  wire  pma_checker_entries_barrier_10_io_x_eff;
  wire  pma_checker_entries_barrier_10_io_x_c;
  wire [19:0] pma_checker_entries_barrier_10_io_y_ppn;
  wire  pma_checker_entries_barrier_10_io_y_u;
  wire  pma_checker_entries_barrier_10_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_10_io_y_ae_final;
  wire  pma_checker_entries_barrier_10_io_y_pf;
  wire  pma_checker_entries_barrier_10_io_y_gf;
  wire  pma_checker_entries_barrier_10_io_y_sw;
  wire  pma_checker_entries_barrier_10_io_y_sx;
  wire  pma_checker_entries_barrier_10_io_y_sr;
  wire  pma_checker_entries_barrier_10_io_y_pw;
  wire  pma_checker_entries_barrier_10_io_y_px;
  wire  pma_checker_entries_barrier_10_io_y_pr;
  wire  pma_checker_entries_barrier_10_io_y_ppp;
  wire  pma_checker_entries_barrier_10_io_y_pal;
  wire  pma_checker_entries_barrier_10_io_y_paa;
  wire  pma_checker_entries_barrier_10_io_y_eff;
  wire  pma_checker_entries_barrier_10_io_y_c;
  wire [19:0] pma_checker_entries_barrier_11_io_x_ppn;
  wire  pma_checker_entries_barrier_11_io_x_u;
  wire  pma_checker_entries_barrier_11_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_11_io_x_ae_final;
  wire  pma_checker_entries_barrier_11_io_x_pf;
  wire  pma_checker_entries_barrier_11_io_x_gf;
  wire  pma_checker_entries_barrier_11_io_x_sw;
  wire  pma_checker_entries_barrier_11_io_x_sx;
  wire  pma_checker_entries_barrier_11_io_x_sr;
  wire  pma_checker_entries_barrier_11_io_x_pw;
  wire  pma_checker_entries_barrier_11_io_x_px;
  wire  pma_checker_entries_barrier_11_io_x_pr;
  wire  pma_checker_entries_barrier_11_io_x_ppp;
  wire  pma_checker_entries_barrier_11_io_x_pal;
  wire  pma_checker_entries_barrier_11_io_x_paa;
  wire  pma_checker_entries_barrier_11_io_x_eff;
  wire  pma_checker_entries_barrier_11_io_x_c;
  wire [19:0] pma_checker_entries_barrier_11_io_y_ppn;
  wire  pma_checker_entries_barrier_11_io_y_u;
  wire  pma_checker_entries_barrier_11_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_11_io_y_ae_final;
  wire  pma_checker_entries_barrier_11_io_y_pf;
  wire  pma_checker_entries_barrier_11_io_y_gf;
  wire  pma_checker_entries_barrier_11_io_y_sw;
  wire  pma_checker_entries_barrier_11_io_y_sx;
  wire  pma_checker_entries_barrier_11_io_y_sr;
  wire  pma_checker_entries_barrier_11_io_y_pw;
  wire  pma_checker_entries_barrier_11_io_y_px;
  wire  pma_checker_entries_barrier_11_io_y_pr;
  wire  pma_checker_entries_barrier_11_io_y_ppp;
  wire  pma_checker_entries_barrier_11_io_y_pal;
  wire  pma_checker_entries_barrier_11_io_y_paa;
  wire  pma_checker_entries_barrier_11_io_y_eff;
  wire  pma_checker_entries_barrier_11_io_y_c;
  wire [19:0] pma_checker_entries_barrier_12_io_x_ppn;
  wire  pma_checker_entries_barrier_12_io_x_u;
  wire  pma_checker_entries_barrier_12_io_x_ae_ptw;
  wire  pma_checker_entries_barrier_12_io_x_ae_final;
  wire  pma_checker_entries_barrier_12_io_x_pf;
  wire  pma_checker_entries_barrier_12_io_x_gf;
  wire  pma_checker_entries_barrier_12_io_x_sw;
  wire  pma_checker_entries_barrier_12_io_x_sx;
  wire  pma_checker_entries_barrier_12_io_x_sr;
  wire  pma_checker_entries_barrier_12_io_x_pw;
  wire  pma_checker_entries_barrier_12_io_x_px;
  wire  pma_checker_entries_barrier_12_io_x_pr;
  wire  pma_checker_entries_barrier_12_io_x_ppp;
  wire  pma_checker_entries_barrier_12_io_x_pal;
  wire  pma_checker_entries_barrier_12_io_x_paa;
  wire  pma_checker_entries_barrier_12_io_x_eff;
  wire  pma_checker_entries_barrier_12_io_x_c;
  wire [19:0] pma_checker_entries_barrier_12_io_y_ppn;
  wire  pma_checker_entries_barrier_12_io_y_u;
  wire  pma_checker_entries_barrier_12_io_y_ae_ptw;
  wire  pma_checker_entries_barrier_12_io_y_ae_final;
  wire  pma_checker_entries_barrier_12_io_y_pf;
  wire  pma_checker_entries_barrier_12_io_y_gf;
  wire  pma_checker_entries_barrier_12_io_y_sw;
  wire  pma_checker_entries_barrier_12_io_y_sx;
  wire  pma_checker_entries_barrier_12_io_y_sr;
  wire  pma_checker_entries_barrier_12_io_y_pw;
  wire  pma_checker_entries_barrier_12_io_y_px;
  wire  pma_checker_entries_barrier_12_io_y_pr;
  wire  pma_checker_entries_barrier_12_io_y_ppp;
  wire  pma_checker_entries_barrier_12_io_y_pal;
  wire  pma_checker_entries_barrier_12_io_y_paa;
  wire  pma_checker_entries_barrier_12_io_y_eff;
  wire  pma_checker_entries_barrier_12_io_y_c;
  wire  lfsr_prng_clock;
  wire  lfsr_prng_reset;
  wire  lfsr_prng_io_increment;
  wire  lfsr_prng_io_out_0;
  wire  lfsr_prng_io_out_1;
  wire  lfsr_prng_io_out_2;
  wire  lfsr_prng_io_out_3;
  wire  lfsr_prng_io_out_4;
  wire  lfsr_prng_io_out_5;
  wire  lfsr_prng_io_out_6;
  wire  lfsr_prng_io_out_7;
  wire  lfsr_prng_io_out_8;
  wire  lfsr_prng_io_out_9;
  wire  lfsr_prng_io_out_10;
  wire  lfsr_prng_io_out_11;
  wire  lfsr_prng_io_out_12;
  wire  lfsr_prng_io_out_13;
  wire  lfsr_prng_io_out_14;
  wire  lfsr_prng_io_out_15;
  wire  metaArb_io_in_0_valid;
  wire [31:0] metaArb_io_in_0_bits_addr;
  wire [5:0] metaArb_io_in_0_bits_idx;
  wire  metaArb_io_in_2_valid;
  wire [31:0] metaArb_io_in_2_bits_addr;
  wire [5:0] metaArb_io_in_2_bits_idx;
  wire [3:0] metaArb_io_in_2_bits_way_en;
  wire [21:0] metaArb_io_in_2_bits_data;
  wire  metaArb_io_in_3_valid;
  wire [31:0] metaArb_io_in_3_bits_addr;
  wire [5:0] metaArb_io_in_3_bits_idx;
  wire [3:0] metaArb_io_in_3_bits_way_en;
  wire [21:0] metaArb_io_in_3_bits_data;
  wire  metaArb_io_in_4_ready;
  wire  metaArb_io_in_4_valid;
  wire [31:0] metaArb_io_in_4_bits_addr;
  wire [5:0] metaArb_io_in_4_bits_idx;
  wire [3:0] metaArb_io_in_4_bits_way_en;
  wire [21:0] metaArb_io_in_4_bits_data;
  wire  metaArb_io_in_5_ready;
  wire  metaArb_io_in_5_valid;
  wire [31:0] metaArb_io_in_5_bits_addr;
  wire [5:0] metaArb_io_in_5_bits_idx;
  wire [3:0] metaArb_io_in_5_bits_way_en;
  wire [21:0] metaArb_io_in_5_bits_data;
  wire  metaArb_io_in_6_ready;
  wire  metaArb_io_in_6_valid;
  wire [31:0] metaArb_io_in_6_bits_addr;
  wire [5:0] metaArb_io_in_6_bits_idx;
  wire [3:0] metaArb_io_in_6_bits_way_en;
  wire [21:0] metaArb_io_in_6_bits_data;
  wire  metaArb_io_in_7_ready;
  wire  metaArb_io_in_7_valid;
  wire [31:0] metaArb_io_in_7_bits_addr;
  wire [5:0] metaArb_io_in_7_bits_idx;
  wire [3:0] metaArb_io_in_7_bits_way_en;
  wire [21:0] metaArb_io_in_7_bits_data;
  wire  metaArb_io_out_valid;
  wire  metaArb_io_out_bits_write;
  wire [31:0] metaArb_io_out_bits_addr;
  wire [5:0] metaArb_io_out_bits_idx;
  wire [3:0] metaArb_io_out_bits_way_en;
  wire [21:0] metaArb_io_out_bits_data;
  wire [31:0] metaArb__GEN_2 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_addr : metaArb_io_in_7_bits_addr;
  wire [5:0] metaArb__GEN_3 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_idx : metaArb_io_in_7_bits_idx;
  wire [3:0] metaArb__GEN_4 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_way_en : metaArb_io_in_7_bits_way_en;
  wire [21:0] metaArb__GEN_5 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_data : metaArb_io_in_7_bits_data;
  wire [31:0] metaArb__GEN_8 = metaArb_io_in_5_valid ? metaArb_io_in_5_bits_addr : metaArb__GEN_2;
  wire [5:0] metaArb__GEN_9 = metaArb_io_in_5_valid ? metaArb_io_in_5_bits_idx : metaArb__GEN_3;
  wire [3:0] metaArb__GEN_10 = metaArb_io_in_5_valid ? metaArb_io_in_5_bits_way_en : metaArb__GEN_4;
  wire [21:0] metaArb__GEN_11 = metaArb_io_in_5_valid ? metaArb_io_in_5_bits_data : metaArb__GEN_5;
  wire [31:0] metaArb__GEN_14 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_addr : metaArb__GEN_8;
  wire [5:0] metaArb__GEN_15 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_idx : metaArb__GEN_9;
  wire [3:0] metaArb__GEN_16 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_way_en : metaArb__GEN_10;
  wire [21:0] metaArb__GEN_17 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_data : metaArb__GEN_11;
  wire  metaArb__GEN_19 = metaArb_io_in_3_valid | metaArb_io_in_4_valid;
  wire [31:0] metaArb__GEN_20 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_addr : metaArb__GEN_14;
  wire [5:0] metaArb__GEN_21 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_idx : metaArb__GEN_15;
  wire [3:0] metaArb__GEN_22 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_way_en : metaArb__GEN_16;
  wire [21:0] metaArb__GEN_23 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_data : metaArb__GEN_17;
  wire  metaArb__GEN_25 = metaArb_io_in_2_valid | metaArb__GEN_19;
  wire [31:0] metaArb__GEN_26 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_addr : metaArb__GEN_20;
  wire [5:0] metaArb__GEN_27 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_idx : metaArb__GEN_21;
  wire [3:0] metaArb__GEN_28 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_way_en : metaArb__GEN_22;
  wire [21:0] metaArb__GEN_29 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_data : metaArb__GEN_23;
  wire  metaArb__grant_T_1 = metaArb_io_in_0_valid | metaArb_io_in_2_valid;
  wire  metaArb__grant_T_2 = metaArb__grant_T_1 | metaArb_io_in_3_valid;
  wire  metaArb__grant_T_3 = metaArb__grant_T_2 | metaArb_io_in_4_valid;
  wire  metaArb__grant_T_4 = metaArb__grant_T_3 | metaArb_io_in_5_valid;
  wire  metaArb__grant_T_5 = metaArb__grant_T_4 | metaArb_io_in_6_valid;
  wire  metaArb_grant_7 = ~metaArb__grant_T_5;
  wire  metaArb__io_out_valid_T = ~metaArb_grant_7;
  wire [5:0] tag_array_RW0_addr;
  wire  tag_array_RW0_en;
  wire  tag_array_RW0_clk;
  wire  tag_array_RW0_wmode;
  wire [21:0] tag_array_RW0_wdata_0;
  wire [21:0] tag_array_RW0_wdata_1;
  wire [21:0] tag_array_RW0_wdata_2;
  wire [21:0] tag_array_RW0_wdata_3;
  wire [21:0] tag_array_RW0_rdata_0;
  wire [21:0] tag_array_RW0_rdata_1;
  wire [21:0] tag_array_RW0_rdata_2;
  wire [21:0] tag_array_RW0_rdata_3;
  wire  tag_array_RW0_wmask_0;
  wire  tag_array_RW0_wmask_1;
  wire  tag_array_RW0_wmask_2;
  wire  tag_array_RW0_wmask_3;
  wire  data_clock;
  wire  data_io_req_valid;
  wire [11:0] data_io_req_bits_addr;
  wire  data_io_req_bits_write;
  wire [31:0] data_io_req_bits_wdata;
  wire [3:0] data_io_req_bits_eccMask;
  wire [3:0] data_io_req_bits_way_en;
  wire [31:0] data_io_resp_0;
  wire [31:0] data_io_resp_1;
  wire [31:0] data_io_resp_2;
  wire [31:0] data_io_resp_3;
  wire  dataArb_io_in_0_valid;
  wire [11:0] dataArb_io_in_0_bits_addr;
  wire  dataArb_io_in_0_bits_write;
  wire [31:0] dataArb_io_in_0_bits_wdata;
  wire [3:0] dataArb_io_in_0_bits_eccMask;
  wire [3:0] dataArb_io_in_0_bits_way_en;
  wire  dataArb_io_in_1_ready;
  wire  dataArb_io_in_1_valid;
  wire [11:0] dataArb_io_in_1_bits_addr;
  wire  dataArb_io_in_1_bits_write;
  wire [31:0] dataArb_io_in_1_bits_wdata;
  wire [3:0] dataArb_io_in_1_bits_way_en;
  wire  dataArb_io_in_2_ready;
  wire  dataArb_io_in_2_valid;
  wire [11:0] dataArb_io_in_2_bits_addr;
  wire [31:0] dataArb_io_in_2_bits_wdata;
  wire  dataArb_io_in_3_ready;
  wire  dataArb_io_in_3_valid;
  wire [11:0] dataArb_io_in_3_bits_addr;
  wire [31:0] dataArb_io_in_3_bits_wdata;
  wire  dataArb_io_out_valid;
  wire [11:0] dataArb_io_out_bits_addr;
  wire  dataArb_io_out_bits_write;
  wire [31:0] dataArb_io_out_bits_wdata;
  wire [3:0] dataArb_io_out_bits_eccMask;
  wire [3:0] dataArb_io_out_bits_way_en;
  wire [11:0] dataArb__GEN_1 = dataArb_io_in_2_valid ? dataArb_io_in_2_bits_addr : dataArb_io_in_3_bits_addr;
  wire [31:0] dataArb__GEN_3 = dataArb_io_in_2_valid ? dataArb_io_in_2_bits_wdata : dataArb_io_in_3_bits_wdata;
  wire [11:0] dataArb__GEN_8 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_addr : dataArb__GEN_1;
  wire  dataArb__GEN_9 = dataArb_io_in_1_valid & dataArb_io_in_1_bits_write;
  wire [31:0] dataArb__GEN_10 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_wdata : dataArb__GEN_3;
  wire [3:0] dataArb__GEN_13 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_way_en : 4'hf;
  wire  dataArb__grant_T = dataArb_io_in_0_valid | dataArb_io_in_1_valid;
  wire  dataArb__grant_T_1 = dataArb__grant_T | dataArb_io_in_2_valid;
  wire  dataArb_grant_3 = ~dataArb__grant_T_1;
  wire  dataArb__io_out_valid_T = ~dataArb_grant_3;
  wire [3:0] amoalu_io_mask;
  wire [4:0] amoalu_io_cmd;
  wire [31:0] amoalu_io_lhs;
  wire [31:0] amoalu_io_rhs;
  wire [31:0] amoalu_io_out;
  wire [7:0] lfsr_lo = {lfsr_prng_io_out_7,lfsr_prng_io_out_6,lfsr_prng_io_out_5,lfsr_prng_io_out_4,lfsr_prng_io_out_3,
    lfsr_prng_io_out_2,lfsr_prng_io_out_1,lfsr_prng_io_out_0};
  wire [15:0] lfsr = {lfsr_prng_io_out_15,lfsr_prng_io_out_14,lfsr_prng_io_out_13,lfsr_prng_io_out_12,
    lfsr_prng_io_out_11,lfsr_prng_io_out_10,lfsr_prng_io_out_9,lfsr_prng_io_out_8,lfsr_lo};
  wire  s1_valid_x12 = io_cpu_req_ready & io_cpu_req_valid;
  reg  s1_valid;
  reg [6:0] lrscCount;
  wire  lrscValid = lrscCount > 7'h3;
  reg  s1_probe;
  reg  s2_probe;
  reg [3:0] release_state;
  wire  releaseInFlight = s1_probe | s2_probe | release_state != 4'h0;
  reg  release_ack_wait;
  reg [31:0] release_ack_addr;
  reg  s2_valid;
  reg [31:0] probe_bits_address;
  wire  s1_valid_masked = s1_valid & ~io_cpu_s1_kill;
  reg [1:0] s2_probe_state_state;
  wire [3:0] _T_138 = {2'h0,s2_probe_state_state};
  wire  _T_195 = 4'h3 == _T_138;
  wire  _T_191 = 4'h2 == _T_138;
  wire  _T_187 = 4'h1 == _T_138;
  wire  _T_183 = 4'h0 == _T_138;
  wire  _T_179 = 4'h7 == _T_138;
  wire  _T_175 = 4'h6 == _T_138;
  wire  _T_171 = 4'h5 == _T_138;
  wire  _T_167 = 4'h4 == _T_138;
  wire  _T_163 = 4'hb == _T_138;
  wire  _T_159 = 4'ha == _T_138;
  wire  _T_155 = 4'h9 == _T_138;
  wire  _T_151 = 4'h8 == _T_138;
  wire  _T_168 = _T_167 ? 1'h0 : _T_163;
  wire  _T_172 = _T_171 ? 1'h0 : _T_168;
  wire  _T_176 = _T_175 ? 1'h0 : _T_172;
  wire  _T_184 = _T_183 ? 1'h0 : _T_179 | _T_176;
  wire  _T_188 = _T_187 ? 1'h0 : _T_184;
  wire  _T_192 = _T_191 ? 1'h0 : _T_188;
  wire  s2_prb_ack_data = _T_195 | _T_192;
  wire  _T_324 = s2_probe_state_state > 2'h0;
  reg [9:0] counter_1;
  wire  _T_329 = release_state == 4'h1;
  wire  _T_330 = release_state == 4'h6;
  wire  _T_331 = release_state == 4'h9;
  wire  _T_333 = _T_329 | _T_330 | _T_331;
  wire [2:0] _GEN_346 = _T_331 ? 3'h6 : 3'h7;
  wire  _T_328 = release_state == 4'h2;
  wire [2:0] _GEN_338 = release_state == 4'h2 ? 3'h5 : 3'h4;
  wire [2:0] tl_out__c_bits_opcode = _T_333 ? _GEN_346 : _GEN_338;
  wire  beats1_opdata_1 = tl_out__c_bits_opcode[0];
  wire [3:0] tl_out__c_bits_size = _T_333 ? 4'h6 : 4'h0;
  wire [26:0] _beats1_decode_T_5 = 27'hfff << tl_out__c_bits_size;
  wire [11:0] _beats1_decode_T_7 = ~_beats1_decode_T_5[11:0];
  wire [9:0] beats1_decode_1 = _beats1_decode_T_7[11:2];
  wire [9:0] beats1_1 = beats1_opdata_1 ? beats1_decode_1 : 10'h0;
  wire  c_last = counter_1 == 10'h1 | beats1_1 == 10'h0;
  reg  s2_release_data_valid;
  wire  c_first = counter_1 == 10'h0;
  wire  _GEN_287 = s2_prb_ack_data ? s2_release_data_valid & ~(c_first & release_ack_wait) : 1'h1;
  wire  _GEN_308 = s2_probe ? _GEN_287 : s2_release_data_valid & ~(c_first & release_ack_wait);
  wire  _GEN_325 = release_state == 4'h5 | _GEN_308;
  wire  tl_out__c_valid = release_state == 4'h3 | _GEN_325;
  wire  _T_318 = auto_out_c_ready & tl_out__c_valid;
  wire  releaseDone = c_last & _T_318;
  wire  _GEN_285 = _T_324 | ~releaseDone;
  wire  probeNack = s2_prb_ack_data | _GEN_285;
  reg [4:0] s1_req_cmd;
  wire  _s1_read_T = s1_req_cmd == 5'h0;
  wire  _s1_read_T_1 = s1_req_cmd == 5'h10;
  wire  _s1_read_T_2 = s1_req_cmd == 5'h6;
  wire  _s1_read_T_3 = s1_req_cmd == 5'h7;
  wire  _s1_read_T_6 = _s1_read_T | _s1_read_T_1 | _s1_read_T_2 | _s1_read_T_3;
  wire  _s1_read_T_7 = s1_req_cmd == 5'h4;
  wire  _s1_read_T_8 = s1_req_cmd == 5'h9;
  wire  _s1_read_T_9 = s1_req_cmd == 5'ha;
  wire  _s1_read_T_10 = s1_req_cmd == 5'hb;
  wire  _s1_read_T_13 = _s1_read_T_7 | _s1_read_T_8 | _s1_read_T_9 | _s1_read_T_10;
  wire  _s1_read_T_14 = s1_req_cmd == 5'h8;
  wire  _s1_read_T_15 = s1_req_cmd == 5'hc;
  wire  _s1_read_T_16 = s1_req_cmd == 5'hd;
  wire  _s1_read_T_17 = s1_req_cmd == 5'he;
  wire  _s1_read_T_18 = s1_req_cmd == 5'hf;
  wire  _s1_read_T_22 = _s1_read_T_14 | _s1_read_T_15 | _s1_read_T_16 | _s1_read_T_17 | _s1_read_T_18;
  wire  _s1_read_T_23 = _s1_read_T_13 | _s1_read_T_22;
  wire  s1_read = _s1_read_T_6 | _s1_read_T_23;
  reg [4:0] s2_req_cmd;
  wire  _s2_write_T_1 = s2_req_cmd == 5'h11;
  wire  _s2_write_T_3 = s2_req_cmd == 5'h7;
  wire  _s2_write_T_5 = s2_req_cmd == 5'h4;
  wire  _s2_write_T_6 = s2_req_cmd == 5'h9;
  wire  _s2_write_T_7 = s2_req_cmd == 5'ha;
  wire  _s2_write_T_8 = s2_req_cmd == 5'hb;
  wire  _s2_write_T_11 = _s2_write_T_5 | _s2_write_T_6 | _s2_write_T_7 | _s2_write_T_8;
  wire  _s2_write_T_12 = s2_req_cmd == 5'h8;
  wire  _s2_write_T_13 = s2_req_cmd == 5'hc;
  wire  _s2_write_T_14 = s2_req_cmd == 5'hd;
  wire  _s2_write_T_15 = s2_req_cmd == 5'he;
  wire  _s2_write_T_16 = s2_req_cmd == 5'hf;
  wire  _s2_write_T_20 = _s2_write_T_12 | _s2_write_T_13 | _s2_write_T_14 | _s2_write_T_15 | _s2_write_T_16;
  wire  _s2_write_T_21 = _s2_write_T_11 | _s2_write_T_20;
  wire  s2_write = s2_req_cmd == 5'h1 | s2_req_cmd == 5'h11 | s2_req_cmd == 5'h7 | _s2_write_T_21;
  reg  pstore1_held;
  wire  pstore1_valid_likely = s2_valid & s2_write | pstore1_held;
  reg [31:0] pstore1_addr;
  reg [31:0] s1_req_addr;
  wire [31:0] s1_vaddr = {s1_req_addr[31:12],s1_req_addr[11:0]};
  wire  _s1_write_T_1 = s1_req_cmd == 5'h11;
  wire  s1_write = s1_req_cmd == 5'h1 | s1_req_cmd == 5'h11 | _s1_read_T_3 | _s1_read_T_23;
  reg [3:0] pstore1_mask;
  wire  _s1_hazard_T_10 = |pstore1_mask[3];
  wire  _s1_hazard_T_9 = |pstore1_mask[2];
  wire  _s1_hazard_T_8 = |pstore1_mask[1];
  wire  _s1_hazard_T_7 = |pstore1_mask[0];
  wire [3:0] _s1_hazard_T_11 = {_s1_hazard_T_10,_s1_hazard_T_9,_s1_hazard_T_8,_s1_hazard_T_7};
  wire [3:0] _s1_hazard_T_16 = {_s1_hazard_T_11[3],_s1_hazard_T_11[2],_s1_hazard_T_11[1],_s1_hazard_T_11[0]};
  reg [1:0] s1_req_size;
  wire  s1_mask_xwr_upper = s1_req_addr[0] | s1_req_size >= 2'h1;
  wire  s1_mask_xwr_lower = s1_req_addr[0] ? 1'h0 : 1'h1;
  wire [1:0] _s1_mask_xwr_T = {s1_mask_xwr_upper,s1_mask_xwr_lower};
  wire [1:0] _s1_mask_xwr_upper_T_5 = s1_req_addr[1] ? _s1_mask_xwr_T : 2'h0;
  wire [1:0] _s1_mask_xwr_upper_T_7 = s1_req_size >= 2'h2 ? 2'h3 : 2'h0;
  wire [1:0] s1_mask_xwr_upper_1 = _s1_mask_xwr_upper_T_5 | _s1_mask_xwr_upper_T_7;
  wire [1:0] s1_mask_xwr_lower_1 = s1_req_addr[1] ? 2'h0 : _s1_mask_xwr_T;
  wire [3:0] s1_mask_xwr = {s1_mask_xwr_upper_1,s1_mask_xwr_lower_1};
  wire  _s1_hazard_T_24 = |s1_mask_xwr[3];
  wire  _s1_hazard_T_23 = |s1_mask_xwr[2];
  wire  _s1_hazard_T_22 = |s1_mask_xwr[1];
  wire  _s1_hazard_T_21 = |s1_mask_xwr[0];
  wire [3:0] _s1_hazard_T_25 = {_s1_hazard_T_24,_s1_hazard_T_23,_s1_hazard_T_22,_s1_hazard_T_21};
  wire [3:0] _s1_hazard_T_30 = {_s1_hazard_T_25[3],_s1_hazard_T_25[2],_s1_hazard_T_25[1],_s1_hazard_T_25[0]};
  wire [3:0] _s1_hazard_T_31 = _s1_hazard_T_16 & _s1_hazard_T_30;
  wire [3:0] _s1_hazard_T_33 = pstore1_mask & s1_mask_xwr;
  wire  _s1_hazard_T_35 = s1_write ? |_s1_hazard_T_31 : |_s1_hazard_T_33;
  wire  _s1_hazard_T_36 = pstore1_addr[11:2] == s1_vaddr[11:2] & _s1_hazard_T_35;
  reg  pstore2_valid;
  reg [31:0] pstore2_addr;
  reg [3:0] mask;
  wire  _s1_hazard_T_48 = |mask[3];
  wire  _s1_hazard_T_47 = |mask[2];
  wire  _s1_hazard_T_46 = |mask[1];
  wire  _s1_hazard_T_45 = |mask[0];
  wire [3:0] _s1_hazard_T_49 = {_s1_hazard_T_48,_s1_hazard_T_47,_s1_hazard_T_46,_s1_hazard_T_45};
  wire [3:0] _s1_hazard_T_54 = {_s1_hazard_T_49[3],_s1_hazard_T_49[2],_s1_hazard_T_49[1],_s1_hazard_T_49[0]};
  wire [3:0] _s1_hazard_T_69 = _s1_hazard_T_54 & _s1_hazard_T_30;
  wire [3:0] _s1_hazard_T_71 = mask & s1_mask_xwr;
  wire  _s1_hazard_T_73 = s1_write ? |_s1_hazard_T_69 : |_s1_hazard_T_71;
  wire  _s1_hazard_T_74 = pstore2_addr[11:2] == s1_vaddr[11:2] & _s1_hazard_T_73;
  wire  _s1_hazard_T_75 = pstore2_valid & _s1_hazard_T_74;
  wire  s1_hazard = pstore1_valid_likely & _s1_hazard_T_36 | _s1_hazard_T_75;
  wire  s1_raw_hazard = s1_read & s1_hazard;
  wire [7:0] _s2_valid_no_xcpt_T = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,
    io_cpu_s2_xcpt_gf_ld,io_cpu_s2_xcpt_gf_st,io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st};
  wire  s2_valid_no_xcpt = s2_valid & ~(|_s2_valid_no_xcpt_T);
  reg  s2_not_nacked_in_s1;
  wire  s2_valid_masked = s2_valid_no_xcpt & s2_not_nacked_in_s1;
  wire  _c_cat_T_48 = s2_req_cmd == 5'h6;
  wire  _c_cat_T_49 = s2_write | s2_req_cmd == 5'h3 | s2_req_cmd == 5'h6;
  reg [1:0] s2_hit_state_state;
  wire [3:0] _T_75 = {s2_write,_c_cat_T_49,s2_hit_state_state};
  wire  _T_133 = 4'h3 == _T_75;
  wire  _T_130 = 4'h2 == _T_75;
  wire  _T_127 = 4'h1 == _T_75;
  wire  _T_124 = 4'h7 == _T_75;
  wire  _T_121 = 4'h6 == _T_75;
  wire  _T_118 = 4'hf == _T_75;
  wire  _T_115 = 4'he == _T_75;
  wire  _T_112 = 4'h0 == _T_75;
  wire  _T_109 = 4'h5 == _T_75;
  wire  _T_106 = 4'h4 == _T_75;
  wire  _T_103 = 4'hd == _T_75;
  wire  _T_100 = 4'hc == _T_75;
  wire  s2_hit = _T_133 | (_T_130 | (_T_127 | (_T_124 | (_T_121 | (_T_118 | _T_115)))));
  wire  s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = s2_valid_masked & s2_hit;
  wire  _s2_read_T = s2_req_cmd == 5'h0;
  wire  _s2_read_T_1 = s2_req_cmd == 5'h10;
  wire  _s2_read_T_6 = _s2_read_T | _s2_read_T_1 | _c_cat_T_48 | _s2_write_T_3;
  wire  s2_read = _s2_read_T_6 | _s2_write_T_21;
  wire  s2_readwrite = s2_read | s2_write;
  wire  s2_valid_hit_pre_data_ecc_and_waw = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_readwrite;
  wire [1:0] _T_102 = _T_100 ? 2'h1 : 2'h0;
  wire [1:0] _T_105 = _T_103 ? 2'h2 : _T_102;
  wire [1:0] _T_108 = _T_106 ? 2'h1 : _T_105;
  wire [1:0] _T_111 = _T_109 ? 2'h2 : _T_108;
  wire [1:0] _T_114 = _T_112 ? 2'h0 : _T_111;
  wire [1:0] _T_117 = _T_115 ? 2'h3 : _T_114;
  wire [1:0] _T_120 = _T_118 ? 2'h3 : _T_117;
  wire [1:0] _T_123 = _T_121 ? 2'h2 : _T_120;
  wire [1:0] _T_126 = _T_124 ? 2'h3 : _T_123;
  wire [1:0] _T_129 = _T_127 ? 2'h1 : _T_126;
  wire [1:0] _T_132 = _T_130 ? 2'h2 : _T_129;
  wire [1:0] s2_grow_param = _T_133 ? 2'h3 : _T_132;
  wire  _s2_update_meta_T = s2_hit_state_state == s2_grow_param;
  wire  s2_update_meta = ~_s2_update_meta_T;
  wire  s1_readwrite = s1_read | s1_write;
  wire  s1_flush_line = s1_req_cmd == 5'h5 & s1_req_size[0];
  wire  s1_cmd_uses_tlb = s1_readwrite | s1_flush_line | s1_req_cmd == 5'h17;
  wire  _T_14 = s1_valid & s1_cmd_uses_tlb & tlb_io_resp_miss;
  wire  _GEN_141 = io_cpu_s2_nack | s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta | _T_14;
  wire  _GEN_161 = s1_valid & s1_raw_hazard | _GEN_141;
  wire  _GEN_306 = probeNack | _GEN_161;
  wire  s1_nack = s2_probe ? _GEN_306 : _GEN_161;
  wire  _s1_valid_not_nacked_T = ~s1_nack;
  wire  s1_valid_not_nacked = s1_valid & ~s1_nack;
  wire  s0_clk_en = metaArb_io_out_valid & ~metaArb_io_out_bits_write;
  wire [31:0] s0_req_addr = {metaArb_io_out_bits_addr[31:6],io_cpu_req_bits_addr[5:0]};
  wire  _T = ~metaArb_io_in_7_ready;
  wire  s0_req_phys = ~metaArb_io_in_7_ready | io_cpu_req_bits_phys;
  reg [6:0] s1_req_tag;
  reg  s1_req_signed;
  reg [1:0] s1_req_dprv;
  reg [31:0] s1_tlb_req_vaddr;
  reg  s1_tlb_req_passthrough;
  reg [1:0] s1_tlb_req_size;
  reg [4:0] s1_tlb_req_cmd;
  reg [1:0] s1_tlb_req_prv;
  wire  s1_sfence = s1_req_cmd == 5'h14 | s1_req_cmd == 5'h15 | s1_req_cmd == 5'h16;
  reg  s1_flush_valid;
  reg  flushed;
  reg  flushing;
  reg [1:0] flushing_req_size;
  reg  cached_grant_wait;
  reg  resetting;
  reg [7:0] flushCounter;
  reg [3:0] refill_way;
  wire  inWriteback = _T_329 | _T_328;
  wire  _io_cpu_req_ready_T = release_state == 4'h0;
  wire  _io_cpu_req_ready_T_1 = ~cached_grant_wait;
  reg  uncachedInFlight_0;
  reg [31:0] uncachedReqs_0_addr;
  reg [6:0] uncachedReqs_0_tag;
  reg [1:0] uncachedReqs_0_size;
  reg  uncachedReqs_0_signed;
  wire  _s0_read_T = io_cpu_req_bits_cmd == 5'h0;
  wire  _s0_read_T_1 = io_cpu_req_bits_cmd == 5'h10;
  wire  _s0_read_T_2 = io_cpu_req_bits_cmd == 5'h6;
  wire  _s0_read_T_3 = io_cpu_req_bits_cmd == 5'h7;
  wire  _s0_read_T_6 = _s0_read_T | _s0_read_T_1 | _s0_read_T_2 | _s0_read_T_3;
  wire  _s0_read_T_7 = io_cpu_req_bits_cmd == 5'h4;
  wire  _s0_read_T_8 = io_cpu_req_bits_cmd == 5'h9;
  wire  _s0_read_T_9 = io_cpu_req_bits_cmd == 5'ha;
  wire  _s0_read_T_10 = io_cpu_req_bits_cmd == 5'hb;
  wire  _s0_read_T_13 = _s0_read_T_7 | _s0_read_T_8 | _s0_read_T_9 | _s0_read_T_10;
  wire  _s0_read_T_14 = io_cpu_req_bits_cmd == 5'h8;
  wire  _s0_read_T_15 = io_cpu_req_bits_cmd == 5'hc;
  wire  _s0_read_T_16 = io_cpu_req_bits_cmd == 5'hd;
  wire  _s0_read_T_17 = io_cpu_req_bits_cmd == 5'he;
  wire  _s0_read_T_18 = io_cpu_req_bits_cmd == 5'hf;
  wire  _s0_read_T_22 = _s0_read_T_14 | _s0_read_T_15 | _s0_read_T_16 | _s0_read_T_17 | _s0_read_T_18;
  wire  _s0_read_T_23 = _s0_read_T_13 | _s0_read_T_22;
  wire  s0_read = _s0_read_T_6 | _s0_read_T_23;
  wire  _dataArb_io_in_3_valid_res_T = io_cpu_req_bits_cmd == 5'h1;
  wire  _dataArb_io_in_3_valid_res_T_1 = io_cpu_req_bits_cmd == 5'h3;
  wire  _dataArb_io_in_3_valid_res_T_2 = _dataArb_io_in_3_valid_res_T | _dataArb_io_in_3_valid_res_T_1;
  wire  res = ~_dataArb_io_in_3_valid_res_T_2;
  wire  _dataArb_io_in_3_valid_T_26 = io_cpu_req_bits_cmd == 5'h11;
  wire  _dataArb_io_in_3_valid_T_47 = _dataArb_io_in_3_valid_res_T | io_cpu_req_bits_cmd == 5'h11 | _s0_read_T_3 |
    _s0_read_T_23;
  wire  _dataArb_io_in_3_valid_T_51 = _dataArb_io_in_3_valid_T_47 & _dataArb_io_in_3_valid_T_26;
  wire  _dataArb_io_in_3_valid_T_52 = s0_read | _dataArb_io_in_3_valid_T_51;
  wire  _dataArb_io_in_3_valid_T_56 = ~reset;
  wire  _dataArb_io_in_3_valid_T_58 = io_cpu_req_valid & res;
  wire [31:0] _dataArb_io_in_3_bits_addr_T_2 = {io_cpu_req_bits_addr[31:12],io_cpu_req_bits_addr[11:0]};
  wire  _GEN_33 = ~dataArb_io_in_3_ready & s0_read ? 1'h0 : release_state == 4'h0 & ~cached_grant_wait &
    _s1_valid_not_nacked_T;
  wire  _s1_did_read_T_54 = dataArb_io_in_3_ready & (io_cpu_req_valid & _dataArb_io_in_3_valid_T_52);
  reg  s1_did_read;
  wire  _GEN_36 = _T ? 1'h0 : _GEN_33;
  wire  _GEN_37 = ~tlb_io_req_ready & ~tlb_io_ptw_resp_valid & ~io_cpu_req_bits_phys ? 1'h0 : _GEN_36;
  wire [31:0] s1_paddr = {tlb_io_resp_paddr[31:12],s1_req_addr[11:0]};
  wire  _T_19 = metaArb_io_out_valid & metaArb_io_out_bits_write;
  wire [21:0] _WIRE_2 = tag_array_RW0_rdata_0;
  wire [19:0] s1_meta_uncorrected_0_tag = _WIRE_2[19:0];
  wire [1:0] s1_meta_uncorrected_0_coh_state = _WIRE_2[21:20];
  wire [21:0] _WIRE_3 = tag_array_RW0_rdata_1;
  wire [19:0] s1_meta_uncorrected_1_tag = _WIRE_3[19:0];
  wire [1:0] s1_meta_uncorrected_1_coh_state = _WIRE_3[21:20];
  wire [21:0] _WIRE_4 = tag_array_RW0_rdata_2;
  wire [19:0] s1_meta_uncorrected_2_tag = _WIRE_4[19:0];
  wire [1:0] s1_meta_uncorrected_2_coh_state = _WIRE_4[21:20];
  wire [21:0] _WIRE_5 = tag_array_RW0_rdata_3;
  wire [19:0] s1_meta_uncorrected_3_tag = _WIRE_5[19:0];
  wire [1:0] s1_meta_uncorrected_3_coh_state = _WIRE_5[21:20];
  wire [19:0] s1_tag = s1_paddr[31:12];
  wire  _T_32 = s1_meta_uncorrected_0_coh_state > 2'h0;
  wire  _T_33 = s1_meta_uncorrected_0_tag == s1_tag;
  wire  _T_34 = _T_32 & s1_meta_uncorrected_0_tag == s1_tag;
  wire  _T_35 = s1_meta_uncorrected_1_coh_state > 2'h0;
  wire  _T_36 = s1_meta_uncorrected_1_tag == s1_tag;
  wire  _T_37 = _T_35 & s1_meta_uncorrected_1_tag == s1_tag;
  wire  _T_38 = s1_meta_uncorrected_2_coh_state > 2'h0;
  wire  _T_39 = s1_meta_uncorrected_2_tag == s1_tag;
  wire  _T_40 = _T_38 & s1_meta_uncorrected_2_tag == s1_tag;
  wire  _T_41 = s1_meta_uncorrected_3_coh_state > 2'h0;
  wire  _T_42 = s1_meta_uncorrected_3_tag == s1_tag;
  wire  _T_43 = _T_41 & s1_meta_uncorrected_3_tag == s1_tag;
  wire [3:0] s1_meta_hit_way = {_T_43,_T_40,_T_37,_T_34};
  wire  _T_45 = ~s1_flush_valid;
  wire [1:0] _T_47 = _T_33 & ~s1_flush_valid ? s1_meta_uncorrected_0_coh_state : 2'h0;
  wire [1:0] _T_51 = _T_36 & ~s1_flush_valid ? s1_meta_uncorrected_1_coh_state : 2'h0;
  wire [1:0] _T_55 = _T_39 & ~s1_flush_valid ? s1_meta_uncorrected_2_coh_state : 2'h0;
  wire [1:0] _T_59 = _T_42 & ~s1_flush_valid ? s1_meta_uncorrected_3_coh_state : 2'h0;
  wire [1:0] _T_60 = _T_47 | _T_51;
  wire [1:0] _T_61 = _T_60 | _T_55;
  wire [1:0] s1_meta_hit_state_state = _T_61 | _T_59;
  wire  s2_hit_valid = s2_hit_state_state > 2'h0;
  reg [3:0] s2_hit_way;
  reg [1:0] s2_victim_way_r;
  wire [3:0] s2_victim_way = 4'h1 << s2_victim_way_r;
  wire [3:0] s2_victim_or_hit_way = s2_hit_valid ? s2_hit_way : s2_victim_way;
  reg [3:0] s2_probe_way;
  wire [3:0] releaseWay = _T_333 ? s2_victim_or_hit_way : s2_probe_way;
  wire [3:0] s1_data_way_x42 = inWriteback ? releaseWay : s1_meta_hit_way;
  wire [15:0] tl_d_data_encoded_lo = {auto_out_d_bits_data[15:8],auto_out_d_bits_data[7:0]};
  wire [15:0] tl_d_data_encoded_hi = {auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16]};
  wire [31:0] _tl_d_data_encoded_T_4 = {auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16],auto_out_d_bits_data[15:
    8],auto_out_d_bits_data[7:0]};
  wire [3:0] _T_67 = ~io_cpu_s1_data_mask;
  wire [3:0] _T_68 = s1_mask_xwr | _T_67;
  wire  s2_valid_x44 = s1_valid_masked & ~s1_sfence;
  reg [31:0] s2_req_addr;
  reg [6:0] s2_req_tag;
  reg [1:0] s2_req_size;
  reg  s2_req_signed;
  reg [1:0] s2_req_dprv;
  wire  _s2_cmd_flush_all_T = s2_req_cmd == 5'h5;
  wire  s2_cmd_flush_all = s2_req_cmd == 5'h5 & ~s2_req_size[0];
  wire  s2_cmd_flush_line = _s2_cmd_flush_all_T & s2_req_size[0];
  reg  s2_tlb_xcpt_pf_ld;
  reg  s2_tlb_xcpt_pf_st;
  reg  s2_tlb_xcpt_ae_ld;
  reg  s2_tlb_xcpt_ae_st;
  reg  s2_tlb_xcpt_ma_ld;
  reg  s2_tlb_xcpt_ma_st;
  reg  s2_pma_cacheable;
  reg [31:0] s2_uncached_resp_addr;
  wire  _T_74 = s1_valid_not_nacked | s1_flush_valid;
  wire [31:0] _GEN_63 = s1_valid_not_nacked | s1_flush_valid ? s1_paddr : s2_req_addr;
  wire [6:0] _GEN_64 = s1_valid_not_nacked | s1_flush_valid ? s1_req_tag : s2_req_tag;
  wire [4:0] _GEN_65 = s1_valid_not_nacked | s1_flush_valid ? s1_req_cmd : s2_req_cmd;
  wire [1:0] _GEN_66 = s1_valid_not_nacked | s1_flush_valid ? s1_req_size : s2_req_size;
  wire  _GEN_67 = s1_valid_not_nacked | s1_flush_valid ? s1_req_signed : s2_req_signed;
  reg [31:0] s2_vaddr_r;
  wire [31:0] s2_vaddr = {s2_vaddr_r[31:12],s2_req_addr[11:0]};
  reg  s2_flush_valid_pre_tag_ecc;
  wire  s1_meta_clk_en = _T_74 | s1_probe;
  reg [21:0] s2_meta_corrected_r;
  wire [19:0] s2_meta_corrected_0_tag = s2_meta_corrected_r[19:0];
  wire [1:0] s2_meta_corrected_0_coh_state = s2_meta_corrected_r[21:20];
  reg [21:0] s2_meta_corrected_r_1;
  wire [19:0] s2_meta_corrected_1_tag = s2_meta_corrected_r_1[19:0];
  wire [1:0] s2_meta_corrected_1_coh_state = s2_meta_corrected_r_1[21:20];
  reg [21:0] s2_meta_corrected_r_2;
  wire [19:0] s2_meta_corrected_2_tag = s2_meta_corrected_r_2[19:0];
  wire [1:0] s2_meta_corrected_2_coh_state = s2_meta_corrected_r_2[21:20];
  reg [21:0] s2_meta_corrected_r_3;
  wire [19:0] s2_meta_corrected_3_tag = s2_meta_corrected_r_3[19:0];
  wire [1:0] s2_meta_corrected_3_coh_state = s2_meta_corrected_r_3[21:20];
  wire  en = s1_valid | inWriteback | io_cpu_replay_next;
  wire  word_en = inWriteback | s1_did_read;
  wire [31:0] s1_all_data_ways_0 = data_io_resp_0;
  wire [31:0] s1_all_data_ways_1 = data_io_resp_1;
  wire [31:0] s1_all_data_ways_2 = data_io_resp_2;
  wire [31:0] s1_all_data_ways_3 = data_io_resp_3;
  wire  s1_word_en = ~io_cpu_replay_next ? word_en : 1'h1;
  wire  grantIsUncachedData = auto_out_d_bits_opcode == 3'h1;
  reg  blockUncachedGrant;
  wire  grantIsRefill = auto_out_d_bits_opcode == 3'h5;
  wire  _T_312 = ~dataArb_io_in_1_ready;
  wire  _grantIsCached_T = auto_out_d_bits_opcode == 3'h4;
  wire  grantIsCached = _grantIsCached_T | grantIsRefill;
  reg [9:0] counter;
  wire  d_first = counter == 10'h0;
  wire  canAcceptCachedGrant = ~_T_333;
  wire  _bundleOut_0_d_ready_T_3 = grantIsCached ? (~d_first | auto_out_e_ready) & canAcceptCachedGrant : 1'h1;
  wire  _GEN_256 = grantIsRefill & ~dataArb_io_in_1_ready ? 1'h0 : _bundleOut_0_d_ready_T_3;
  wire  tl_out__d_ready = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? 1'h0 : _GEN_256;
  wire  _T_292 = tl_out__d_ready & auto_out_d_valid;
  wire  _T_288 = auto_out_d_bits_opcode == 3'h0;
  wire  _T_289 = auto_out_d_bits_opcode == 3'h2;
  wire  grantIsUncached = grantIsUncachedData | _T_288 | _T_289;
  wire [4:0] _GEN_212 = grantIsUncachedData ? 5'h10 : {{1'd0}, s1_data_way_x42};
  wire [4:0] _GEN_221 = grantIsUncached ? _GEN_212 : {{1'd0}, s1_data_way_x42};
  wire [4:0] _GEN_234 = grantIsCached ? {{1'd0}, s1_data_way_x42} : _GEN_221;
  wire [4:0] s1_data_way = _T_292 ? _GEN_234 : {{1'd0}, s1_data_way_x42};
  wire [4:0] _s2_data_T_1 = s1_word_en ? s1_data_way : 5'h0;
  wire [31:0] _s2_data_T_7 = _s2_data_T_1[0] ? s1_all_data_ways_0 : 32'h0;
  wire [31:0] _s2_data_T_8 = _s2_data_T_1[1] ? s1_all_data_ways_1 : 32'h0;
  wire [31:0] _s2_data_T_9 = _s2_data_T_1[2] ? s1_all_data_ways_2 : 32'h0;
  wire [31:0] _s2_data_T_10 = _s2_data_T_1[3] ? s1_all_data_ways_3 : 32'h0;
  wire [31:0] _s2_data_T_11 = _s2_data_T_1[4] ? _tl_d_data_encoded_T_4 : 32'h0;
  wire [31:0] _s2_data_T_12 = _s2_data_T_7 | _s2_data_T_8;
  wire [31:0] _s2_data_T_13 = _s2_data_T_12 | _s2_data_T_9;
  wire [31:0] _s2_data_T_14 = _s2_data_T_13 | _s2_data_T_10;
  wire [31:0] _s2_data_T_15 = _s2_data_T_14 | _s2_data_T_11;
  reg [31:0] s2_data;
  wire [15:0] s2_data_corrected_lo = {s2_data[15:8],s2_data[7:0]};
  wire [15:0] s2_data_corrected_hi = {s2_data[31:24],s2_data[23:16]};
  wire [31:0] s2_data_corrected = {s2_data[31:24],s2_data[23:16],s2_data[15:8],s2_data[7:0]};
  wire  s2_valid_flush_line = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_cmd_flush_line;
  wire  _s2_valid_miss_T_3 = ~s2_hit;
  wire  s2_valid_miss = s2_valid_masked & s2_readwrite & ~s2_hit;
  wire  s2_uncached = ~s2_pma_cacheable;
  wire  _s2_valid_cached_miss_T = ~s2_uncached;
  wire  _s2_valid_cached_miss_T_2 = |uncachedInFlight_0;
  wire  _s2_valid_cached_miss_T_3 = ~(|uncachedInFlight_0);
  wire  s2_valid_cached_miss = s2_valid_miss & ~s2_uncached & ~(|uncachedInFlight_0);
  wire  s2_want_victimize = s2_valid_cached_miss | s2_valid_flush_line | s2_flush_valid_pre_tag_ecc;
  wire  _s2_cannot_victimize_T = ~s2_flush_valid_pre_tag_ecc;
  wire  s2_valid_uncached_pending = s2_valid_miss & s2_uncached & ~(&uncachedInFlight_0);
  wire [19:0] _s2_victim_tag_T_6 = s2_victim_way[0] ? s2_meta_corrected_0_tag : 20'h0;
  wire [19:0] _s2_victim_tag_T_7 = s2_victim_way[1] ? s2_meta_corrected_1_tag : 20'h0;
  wire [19:0] _s2_victim_tag_T_8 = s2_victim_way[2] ? s2_meta_corrected_2_tag : 20'h0;
  wire [19:0] _s2_victim_tag_T_9 = s2_victim_way[3] ? s2_meta_corrected_3_tag : 20'h0;
  wire [19:0] _s2_victim_tag_T_10 = _s2_victim_tag_T_6 | _s2_victim_tag_T_7;
  wire [19:0] _s2_victim_tag_T_11 = _s2_victim_tag_T_10 | _s2_victim_tag_T_8;
  wire [19:0] _s2_victim_tag_T_12 = _s2_victim_tag_T_11 | _s2_victim_tag_T_9;
  wire [1:0] _s2_victim_tag_T_13 = s2_victim_way[0] ? s2_meta_corrected_0_coh_state : 2'h0;
  wire [1:0] _s2_victim_tag_T_14 = s2_victim_way[1] ? s2_meta_corrected_1_coh_state : 2'h0;
  wire [1:0] _s2_victim_tag_T_15 = s2_victim_way[2] ? s2_meta_corrected_2_coh_state : 2'h0;
  wire [1:0] _s2_victim_tag_T_16 = s2_victim_way[3] ? s2_meta_corrected_3_coh_state : 2'h0;
  wire [1:0] _s2_victim_tag_T_17 = _s2_victim_tag_T_13 | _s2_victim_tag_T_14;
  wire [1:0] _s2_victim_tag_T_18 = _s2_victim_tag_T_17 | _s2_victim_tag_T_15;
  wire [1:0] _s2_victim_tag_T_19 = _s2_victim_tag_T_18 | _s2_victim_tag_T_16;
  wire [19:0] s2_victim_tag = s2_valid_flush_line ? s2_req_addr[31:12] : _s2_victim_tag_T_12;
  wire [1:0] s2_victim_state_state = s2_hit_valid ? s2_hit_state_state : _s2_victim_tag_T_19;
  wire [2:0] _T_153 = _T_151 ? 3'h5 : 3'h0;
  wire [2:0] _T_157 = _T_155 ? 3'h2 : _T_153;
  wire [2:0] _T_161 = _T_159 ? 3'h1 : _T_157;
  wire [2:0] _T_165 = _T_163 ? 3'h1 : _T_161;
  wire [2:0] _T_169 = _T_167 ? 3'h5 : _T_165;
  wire [2:0] _T_173 = _T_171 ? 3'h4 : _T_169;
  wire [1:0] _T_174 = _T_171 ? 2'h1 : 2'h0;
  wire [2:0] _T_177 = _T_175 ? 3'h0 : _T_173;
  wire [1:0] _T_178 = _T_175 ? 2'h1 : _T_174;
  wire [2:0] _T_181 = _T_179 ? 3'h0 : _T_177;
  wire [1:0] _T_182 = _T_179 ? 2'h1 : _T_178;
  wire [2:0] _T_185 = _T_183 ? 3'h5 : _T_181;
  wire [1:0] _T_186 = _T_183 ? 2'h0 : _T_182;
  wire [2:0] _T_189 = _T_187 ? 3'h4 : _T_185;
  wire [1:0] _T_190 = _T_187 ? 2'h1 : _T_186;
  wire [2:0] _T_193 = _T_191 ? 3'h3 : _T_189;
  wire [1:0] _T_194 = _T_191 ? 2'h2 : _T_190;
  wire [2:0] s2_report_param = _T_195 ? 3'h3 : _T_193;
  wire [1:0] probeNewCoh_state = _T_195 ? 2'h2 : _T_194;
  wire [3:0] _T_203 = {2'h2,s2_victim_state_state};
  wire  _T_216 = 4'h8 == _T_203;
  wire [2:0] _T_218 = _T_216 ? 3'h5 : 3'h0;
  wire  _T_220 = 4'h9 == _T_203;
  wire [2:0] _T_222 = _T_220 ? 3'h2 : _T_218;
  wire  _T_224 = 4'ha == _T_203;
  wire [2:0] _T_226 = _T_224 ? 3'h1 : _T_222;
  wire  _T_228 = 4'hb == _T_203;
  wire [2:0] _T_230 = _T_228 ? 3'h1 : _T_226;
  wire  _T_232 = 4'h4 == _T_203;
  wire  _T_233 = _T_232 ? 1'h0 : _T_228;
  wire [2:0] _T_234 = _T_232 ? 3'h5 : _T_230;
  wire  _T_236 = 4'h5 == _T_203;
  wire  _T_237 = _T_236 ? 1'h0 : _T_233;
  wire [2:0] _T_238 = _T_236 ? 3'h4 : _T_234;
  wire [1:0] _T_239 = _T_236 ? 2'h1 : 2'h0;
  wire  _T_240 = 4'h6 == _T_203;
  wire  _T_241 = _T_240 ? 1'h0 : _T_237;
  wire [2:0] _T_242 = _T_240 ? 3'h0 : _T_238;
  wire [1:0] _T_243 = _T_240 ? 2'h1 : _T_239;
  wire  _T_244 = 4'h7 == _T_203;
  wire [2:0] _T_246 = _T_244 ? 3'h0 : _T_242;
  wire [1:0] _T_247 = _T_244 ? 2'h1 : _T_243;
  wire  _T_248 = 4'h0 == _T_203;
  wire  _T_249 = _T_248 ? 1'h0 : _T_244 | _T_241;
  wire [2:0] _T_250 = _T_248 ? 3'h5 : _T_246;
  wire [1:0] _T_251 = _T_248 ? 2'h0 : _T_247;
  wire  _T_252 = 4'h1 == _T_203;
  wire  _T_253 = _T_252 ? 1'h0 : _T_249;
  wire [2:0] _T_254 = _T_252 ? 3'h4 : _T_250;
  wire [1:0] _T_255 = _T_252 ? 2'h1 : _T_251;
  wire  _T_256 = 4'h2 == _T_203;
  wire  _T_257 = _T_256 ? 1'h0 : _T_253;
  wire [2:0] _T_258 = _T_256 ? 3'h3 : _T_254;
  wire [1:0] _T_259 = _T_256 ? 2'h2 : _T_255;
  wire  _T_260 = 4'h3 == _T_203;
  wire  s2_victim_dirty = _T_260 | _T_257;
  wire [2:0] s2_shrink_param = _T_260 ? 3'h3 : _T_258;
  wire [1:0] voluntaryNewCoh_state = _T_260 ? 2'h2 : _T_259;
  wire  s2_dont_nack_uncached = s2_valid_uncached_pending & auto_out_a_ready;
  wire  _s2_dont_nack_misc_T_8 = s2_cmd_flush_line & _s2_valid_miss_T_3;
  wire  _s2_dont_nack_misc_T_9 = s2_cmd_flush_all & flushed & ~flushing | _s2_dont_nack_misc_T_8;
  wire  _s2_dont_nack_misc_T_10 = s2_req_cmd == 5'h17;
  wire  _s2_dont_nack_misc_T_11 = _s2_dont_nack_misc_T_9 | _s2_dont_nack_misc_T_10;
  wire  s2_dont_nack_misc = s2_valid_masked & _s2_dont_nack_misc_T_11;
  wire  _io_cpu_s2_nack_T_4 = ~s2_valid_hit_pre_data_ecc_and_waw;
  wire [19:0] metaArb_io_in_2_bits_data_meta_tag = s2_req_addr[31:12];
  wire  _lrscBackingOff_T = lrscCount > 7'h0;
  reg [25:0] lrscAddr;
  wire  lrscAddrMatch = lrscAddr == s2_req_addr[31:6];
  wire  s2_sc_fail = _s2_write_T_3 & ~(lrscValid & lrscAddrMatch);
  wire [6:0] _lrscCount_T = s2_hit ? 7'h4f : 7'h0;
  wire [6:0] _GEN_143 = s2_valid_hit_pre_data_ecc_and_waw & _c_cat_T_48 & _io_cpu_req_ready_T_1 | s2_valid_cached_miss
     ? _lrscCount_T : lrscCount;
  wire [6:0] _lrscCount_T_2 = lrscCount - 7'h1;
  wire  _pstore1_cmd_T = s1_valid_not_nacked & s1_write;
  reg [4:0] pstore1_cmd;
  reg [31:0] pstore1_data;
  reg [3:0] pstore1_way;
  wire  _pstore1_rmw_T_51 = s1_write & _s1_write_T_1;
  wire  _pstore1_rmw_T_52 = s1_read | _pstore1_rmw_T_51;
  reg  pstore1_rmw_r;
  wire  _pstore1_merge_T = s2_valid_hit_pre_data_ecc_and_waw & s2_write;
  wire  _pstore1_merge_T_2 = s2_valid_hit_pre_data_ecc_and_waw & s2_write & ~s2_sc_fail;
  wire  pstore_drain_opportunistic = ~_dataArb_io_in_3_valid_T_58;
  reg  pstore_drain_on_miss_REG;
  wire  pstore_drain_on_miss = releaseInFlight | pstore_drain_on_miss_REG;
  wire  pstore1_valid = _pstore1_merge_T_2 | pstore1_held;
  wire  pstore_drain_structural = pstore1_valid_likely & pstore2_valid & (s1_valid & s1_write | pstore1_rmw_r);
  wire  _T_275 = _pstore1_merge_T | pstore1_held;
  wire  _pstore_drain_T_10 = (_T_275 & ~pstore1_rmw_r | pstore2_valid) & (pstore_drain_opportunistic |
    pstore_drain_on_miss);
  wire  pstore_drain = pstore_drain_structural | _pstore_drain_T_10;
  wire  _pstore1_held_T_9 = ~pstore_drain;
  wire  advance_pstore1 = pstore1_valid & pstore2_valid == pstore_drain;
  reg [3:0] pstore2_way;
  wire [31:0] pstore1_storegen_data = amoalu_io_out;
  reg [7:0] pstore2_storegen_data_r;
  reg [7:0] pstore2_storegen_data_r_1;
  reg [7:0] pstore2_storegen_data_r_2;
  reg [7:0] pstore2_storegen_data_r_3;
  wire [31:0] pstore2_storegen_data = {pstore2_storegen_data_r_3,pstore2_storegen_data_r_2,pstore2_storegen_data_r_1,
    pstore2_storegen_data_r};
  wire [3:0] _pstore2_storegen_mask_mask_T = ~pstore1_mask;
  wire [3:0] _pstore2_storegen_mask_mask_T_2 = ~_pstore2_storegen_mask_mask_T;
  wire [31:0] _dataArb_io_in_0_bits_addr_T = pstore2_valid ? pstore2_addr : pstore1_addr;
  wire [31:0] _dataArb_io_in_0_bits_wdata_T = pstore2_valid ? pstore2_storegen_data : pstore1_data;
  wire [15:0] dataArb_io_in_0_bits_wdata_lo = {_dataArb_io_in_0_bits_wdata_T[15:8],_dataArb_io_in_0_bits_wdata_T[7:0]};
  wire [15:0] dataArb_io_in_0_bits_wdata_hi = {_dataArb_io_in_0_bits_wdata_T[31:24],_dataArb_io_in_0_bits_wdata_T[23:16]
    };
  wire [3:0] _dataArb_io_in_0_bits_eccMask_T = pstore2_valid ? mask : pstore1_mask;
  wire  _dataArb_io_in_0_bits_eccMask_T_5 = |_dataArb_io_in_0_bits_eccMask_T[0];
  wire  _dataArb_io_in_0_bits_eccMask_T_6 = |_dataArb_io_in_0_bits_eccMask_T[1];
  wire  _dataArb_io_in_0_bits_eccMask_T_7 = |_dataArb_io_in_0_bits_eccMask_T[2];
  wire  _dataArb_io_in_0_bits_eccMask_T_8 = |_dataArb_io_in_0_bits_eccMask_T[3];
  wire [1:0] dataArb_io_in_0_bits_eccMask_lo = {_dataArb_io_in_0_bits_eccMask_T_6,_dataArb_io_in_0_bits_eccMask_T_5};
  wire [1:0] dataArb_io_in_0_bits_eccMask_hi = {_dataArb_io_in_0_bits_eccMask_T_8,_dataArb_io_in_0_bits_eccMask_T_7};
  wire  _a_source_T = ~uncachedInFlight_0;
  wire [1:0] _a_source_T_1 = {_a_source_T, 1'h0};
  wire  a_source = _a_source_T_1[0] ? 1'h0 : 1'h1;
  wire [31:0] acquire_address = {s2_req_addr[31:6], 6'h0};
  wire [18:0] a_mask = {{15'd0}, pstore1_mask};
  wire [1:0] _get_a_mask_sizeOH_T_1 = 2'h1 << s2_req_size[0];
  wire [1:0] get_a_mask_sizeOH = _get_a_mask_sizeOH_T_1 | 2'h1;
  wire  _get_a_mask_T = s2_req_size >= 2'h2;
  wire  get_a_mask_size = get_a_mask_sizeOH[1];
  wire  get_a_mask_bit = s2_req_addr[1];
  wire  get_a_mask_nbit = ~get_a_mask_bit;
  wire  get_a_mask_acc = _get_a_mask_T | get_a_mask_size & get_a_mask_nbit;
  wire  get_a_mask_acc_1 = _get_a_mask_T | get_a_mask_size & get_a_mask_bit;
  wire  get_a_mask_size_1 = get_a_mask_sizeOH[0];
  wire  get_a_mask_bit_1 = s2_req_addr[0];
  wire  get_a_mask_nbit_1 = ~get_a_mask_bit_1;
  wire  get_a_mask_eq_2 = get_a_mask_nbit & get_a_mask_nbit_1;
  wire  get_a_mask_acc_2 = get_a_mask_acc | get_a_mask_size_1 & get_a_mask_eq_2;
  wire  get_a_mask_eq_3 = get_a_mask_nbit & get_a_mask_bit_1;
  wire  get_a_mask_acc_3 = get_a_mask_acc | get_a_mask_size_1 & get_a_mask_eq_3;
  wire  get_a_mask_eq_4 = get_a_mask_bit & get_a_mask_nbit_1;
  wire  get_a_mask_acc_4 = get_a_mask_acc_1 | get_a_mask_size_1 & get_a_mask_eq_4;
  wire  get_a_mask_eq_5 = get_a_mask_bit & get_a_mask_bit_1;
  wire  get_a_mask_acc_5 = get_a_mask_acc_1 | get_a_mask_size_1 & get_a_mask_eq_5;
  wire [3:0] get_mask = {get_a_mask_acc_5,get_a_mask_acc_4,get_a_mask_acc_3,get_a_mask_acc_2};
  wire [2:0] _atomics_T_1_opcode = 5'h4 == s2_req_cmd ? 3'h3 : 3'h0;
  wire [3:0] atomics_a_size = {{2'd0}, s2_req_size};
  wire [3:0] _atomics_T_1_size = 5'h4 == s2_req_cmd ? atomics_a_size : 4'h0;
  wire [31:0] _atomics_T_1_address = 5'h4 == s2_req_cmd ? s2_req_addr : 32'h0;
  wire [3:0] _atomics_T_1_mask = 5'h4 == s2_req_cmd ? get_mask : 4'h0;
  wire [31:0] _atomics_T_1_data = 5'h4 == s2_req_cmd ? pstore1_data : 32'h0;
  wire [2:0] _atomics_T_3_opcode = 5'h9 == s2_req_cmd ? 3'h3 : _atomics_T_1_opcode;
  wire [2:0] _atomics_T_3_param = 5'h9 == s2_req_cmd ? 3'h0 : _atomics_T_1_opcode;
  wire [3:0] _atomics_T_3_size = 5'h9 == s2_req_cmd ? atomics_a_size : _atomics_T_1_size;
  wire  _atomics_T_3_source = 5'h9 == s2_req_cmd ? a_source : 5'h4 == s2_req_cmd & a_source;
  wire [31:0] _atomics_T_3_address = 5'h9 == s2_req_cmd ? s2_req_addr : _atomics_T_1_address;
  wire [3:0] _atomics_T_3_mask = 5'h9 == s2_req_cmd ? get_mask : _atomics_T_1_mask;
  wire [31:0] _atomics_T_3_data = 5'h9 == s2_req_cmd ? pstore1_data : _atomics_T_1_data;
  wire [2:0] _atomics_T_5_opcode = 5'ha == s2_req_cmd ? 3'h3 : _atomics_T_3_opcode;
  wire [2:0] _atomics_T_5_param = 5'ha == s2_req_cmd ? 3'h1 : _atomics_T_3_param;
  wire [3:0] _atomics_T_5_size = 5'ha == s2_req_cmd ? atomics_a_size : _atomics_T_3_size;
  wire  _atomics_T_5_source = 5'ha == s2_req_cmd ? a_source : _atomics_T_3_source;
  wire [31:0] _atomics_T_5_address = 5'ha == s2_req_cmd ? s2_req_addr : _atomics_T_3_address;
  wire [3:0] _atomics_T_5_mask = 5'ha == s2_req_cmd ? get_mask : _atomics_T_3_mask;
  wire [31:0] _atomics_T_5_data = 5'ha == s2_req_cmd ? pstore1_data : _atomics_T_3_data;
  wire [2:0] _atomics_T_7_opcode = 5'hb == s2_req_cmd ? 3'h3 : _atomics_T_5_opcode;
  wire [2:0] _atomics_T_7_param = 5'hb == s2_req_cmd ? 3'h2 : _atomics_T_5_param;
  wire [3:0] _atomics_T_7_size = 5'hb == s2_req_cmd ? atomics_a_size : _atomics_T_5_size;
  wire  _atomics_T_7_source = 5'hb == s2_req_cmd ? a_source : _atomics_T_5_source;
  wire [31:0] _atomics_T_7_address = 5'hb == s2_req_cmd ? s2_req_addr : _atomics_T_5_address;
  wire [3:0] _atomics_T_7_mask = 5'hb == s2_req_cmd ? get_mask : _atomics_T_5_mask;
  wire [31:0] _atomics_T_7_data = 5'hb == s2_req_cmd ? pstore1_data : _atomics_T_5_data;
  wire [2:0] _atomics_T_9_opcode = 5'h8 == s2_req_cmd ? 3'h2 : _atomics_T_7_opcode;
  wire [2:0] _atomics_T_9_param = 5'h8 == s2_req_cmd ? 3'h4 : _atomics_T_7_param;
  wire [3:0] _atomics_T_9_size = 5'h8 == s2_req_cmd ? atomics_a_size : _atomics_T_7_size;
  wire  _atomics_T_9_source = 5'h8 == s2_req_cmd ? a_source : _atomics_T_7_source;
  wire [31:0] _atomics_T_9_address = 5'h8 == s2_req_cmd ? s2_req_addr : _atomics_T_7_address;
  wire [3:0] _atomics_T_9_mask = 5'h8 == s2_req_cmd ? get_mask : _atomics_T_7_mask;
  wire [31:0] _atomics_T_9_data = 5'h8 == s2_req_cmd ? pstore1_data : _atomics_T_7_data;
  wire [2:0] _atomics_T_11_opcode = 5'hc == s2_req_cmd ? 3'h2 : _atomics_T_9_opcode;
  wire [2:0] _atomics_T_11_param = 5'hc == s2_req_cmd ? 3'h0 : _atomics_T_9_param;
  wire [3:0] _atomics_T_11_size = 5'hc == s2_req_cmd ? atomics_a_size : _atomics_T_9_size;
  wire  _atomics_T_11_source = 5'hc == s2_req_cmd ? a_source : _atomics_T_9_source;
  wire [31:0] _atomics_T_11_address = 5'hc == s2_req_cmd ? s2_req_addr : _atomics_T_9_address;
  wire [3:0] _atomics_T_11_mask = 5'hc == s2_req_cmd ? get_mask : _atomics_T_9_mask;
  wire [31:0] _atomics_T_11_data = 5'hc == s2_req_cmd ? pstore1_data : _atomics_T_9_data;
  wire [2:0] _atomics_T_13_opcode = 5'hd == s2_req_cmd ? 3'h2 : _atomics_T_11_opcode;
  wire [2:0] _atomics_T_13_param = 5'hd == s2_req_cmd ? 3'h1 : _atomics_T_11_param;
  wire [3:0] _atomics_T_13_size = 5'hd == s2_req_cmd ? atomics_a_size : _atomics_T_11_size;
  wire  _atomics_T_13_source = 5'hd == s2_req_cmd ? a_source : _atomics_T_11_source;
  wire [31:0] _atomics_T_13_address = 5'hd == s2_req_cmd ? s2_req_addr : _atomics_T_11_address;
  wire [3:0] _atomics_T_13_mask = 5'hd == s2_req_cmd ? get_mask : _atomics_T_11_mask;
  wire [31:0] _atomics_T_13_data = 5'hd == s2_req_cmd ? pstore1_data : _atomics_T_11_data;
  wire [2:0] _atomics_T_15_opcode = 5'he == s2_req_cmd ? 3'h2 : _atomics_T_13_opcode;
  wire [2:0] _atomics_T_15_param = 5'he == s2_req_cmd ? 3'h2 : _atomics_T_13_param;
  wire [3:0] _atomics_T_15_size = 5'he == s2_req_cmd ? atomics_a_size : _atomics_T_13_size;
  wire  _atomics_T_15_source = 5'he == s2_req_cmd ? a_source : _atomics_T_13_source;
  wire [31:0] _atomics_T_15_address = 5'he == s2_req_cmd ? s2_req_addr : _atomics_T_13_address;
  wire [3:0] _atomics_T_15_mask = 5'he == s2_req_cmd ? get_mask : _atomics_T_13_mask;
  wire [31:0] _atomics_T_15_data = 5'he == s2_req_cmd ? pstore1_data : _atomics_T_13_data;
  wire [2:0] atomics_opcode = 5'hf == s2_req_cmd ? 3'h2 : _atomics_T_15_opcode;
  wire [2:0] atomics_param = 5'hf == s2_req_cmd ? 3'h3 : _atomics_T_15_param;
  wire [3:0] atomics_size = 5'hf == s2_req_cmd ? atomics_a_size : _atomics_T_15_size;
  wire  atomics_source = 5'hf == s2_req_cmd ? a_source : _atomics_T_15_source;
  wire [31:0] atomics_address = 5'hf == s2_req_cmd ? s2_req_addr : _atomics_T_15_address;
  wire [3:0] atomics_mask = 5'hf == s2_req_cmd ? get_mask : _atomics_T_15_mask;
  wire [31:0] atomics_data = 5'hf == s2_req_cmd ? pstore1_data : _atomics_T_15_data;
  wire [31:0] _tl_out_a_valid_T_1 = s2_req_addr ^ release_ack_addr;
  wire  _tl_out_a_valid_T_5 = ~(release_ack_wait & _tl_out_a_valid_T_1[21:6] == 16'h0);
  wire  _tl_out_a_valid_T_6 = s2_valid_cached_miss & _tl_out_a_valid_T_5;
  wire  _tl_out_a_valid_T_7 = ~release_ack_wait;
  wire  _tl_out_a_valid_T_10 = ~s2_victim_dirty;
  wire  _tl_out_a_valid_T_12 = _tl_out_a_valid_T_6 & _tl_out_a_valid_T_10;
  wire  tl_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12;
  wire [2:0] _tl_out_a_bits_T_6_opcode = ~s2_read ? 3'h0 : atomics_opcode;
  wire [2:0] _tl_out_a_bits_T_6_param = ~s2_read ? 3'h0 : atomics_param;
  wire [3:0] _tl_out_a_bits_T_6_size = ~s2_read ? atomics_a_size : atomics_size;
  wire  _tl_out_a_bits_T_6_source = ~s2_read ? a_source : atomics_source;
  wire [31:0] _tl_out_a_bits_T_6_address = ~s2_read ? s2_req_addr : atomics_address;
  wire [3:0] _tl_out_a_bits_T_6_mask = ~s2_read ? get_mask : atomics_mask;
  wire [31:0] _tl_out_a_bits_T_6_data = ~s2_read ? pstore1_data : atomics_data;
  wire [2:0] _tl_out_a_bits_T_7_opcode = _s2_write_T_1 ? 3'h1 : _tl_out_a_bits_T_6_opcode;
  wire [2:0] _tl_out_a_bits_T_7_param = _s2_write_T_1 ? 3'h0 : _tl_out_a_bits_T_6_param;
  wire [3:0] _tl_out_a_bits_T_7_size = _s2_write_T_1 ? atomics_a_size : _tl_out_a_bits_T_6_size;
  wire  _tl_out_a_bits_T_7_source = _s2_write_T_1 ? a_source : _tl_out_a_bits_T_6_source;
  wire [31:0] _tl_out_a_bits_T_7_address = _s2_write_T_1 ? s2_req_addr : _tl_out_a_bits_T_6_address;
  wire [3:0] putpartial_mask = a_mask[3:0];
  wire [3:0] _tl_out_a_bits_T_7_mask = _s2_write_T_1 ? putpartial_mask : _tl_out_a_bits_T_6_mask;
  wire [31:0] _tl_out_a_bits_T_7_data = _s2_write_T_1 ? pstore1_data : _tl_out_a_bits_T_6_data;
  wire [2:0] _tl_out_a_bits_T_8_opcode = ~s2_write ? 3'h4 : _tl_out_a_bits_T_7_opcode;
  wire [2:0] _tl_out_a_bits_T_8_param = ~s2_write ? 3'h0 : _tl_out_a_bits_T_7_param;
  wire [3:0] _tl_out_a_bits_T_8_size = ~s2_write ? atomics_a_size : _tl_out_a_bits_T_7_size;
  wire  _tl_out_a_bits_T_8_source = ~s2_write ? a_source : _tl_out_a_bits_T_7_source;
  wire [31:0] _tl_out_a_bits_T_8_address = ~s2_write ? s2_req_addr : _tl_out_a_bits_T_7_address;
  wire [3:0] _tl_out_a_bits_T_8_mask = ~s2_write ? get_mask : _tl_out_a_bits_T_7_mask;
  wire [31:0] _tl_out_a_bits_T_8_data = ~s2_write ? 32'h0 : _tl_out_a_bits_T_7_data;
  wire [2:0] tl_out_a_bits_a_param = {{1'd0}, s2_grow_param};
  wire [1:0] _a_sel_T = 2'h1 << a_source;
  wire  a_sel = _a_sel_T[1];
  wire  _T_284 = auto_out_a_ready & tl_out_a_valid;
  wire  _GEN_162 = a_sel | uncachedInFlight_0;
  wire  _GEN_175 = s2_uncached ? _GEN_162 : uncachedInFlight_0;
  wire  _GEN_188 = s2_uncached ? cached_grant_wait : 1'h1;
  wire  _GEN_190 = _T_284 ? _GEN_175 : uncachedInFlight_0;
  wire  _GEN_203 = _T_284 ? _GEN_188 : cached_grant_wait;
  wire [26:0] _beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size;
  wire [11:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[11:0];
  wire [9:0] beats1_decode = _beats1_decode_T_3[11:2];
  wire  beats1_opdata = auto_out_d_bits_opcode[0];
  wire [9:0] beats1 = beats1_opdata ? beats1_decode : 10'h0;
  wire [9:0] counter1 = counter - 10'h1;
  wire  d_last = counter == 10'h1 | beats1 == 10'h0;
  wire  d_done = d_last & _T_292;
  wire [9:0] _count_T = ~counter1;
  wire [9:0] count = beats1 & _count_T;
  wire [11:0] d_address_inc = {count, 2'h0};
  wire  _tl_d_data_encoded_T_8 = ~grantIsUncached;
  wire  grantIsVoluntary = auto_out_d_bits_opcode == 3'h6;
  wire [1:0] _uncachedRespIdxOH_T = 2'h1 << auto_out_d_bits_source;
  wire  uncachedRespIdxOH = _uncachedRespIdxOH_T[1];
  wire  _T_297 = uncachedRespIdxOH & d_last;
  wire  _GEN_211 = uncachedRespIdxOH & d_last ? 1'h0 : _GEN_190;
  wire [31:0] dontCareBits = {s1_paddr[31:2], 2'h0};
  wire [31:0] _GEN_451 = {{30'd0}, uncachedReqs_0_addr[1:0]};
  wire [31:0] _s2_req_addr_T_1 = dontCareBits | _GEN_451;
  wire  _GEN_219 = grantIsVoluntary ? 1'h0 : release_ack_wait;
  wire  _GEN_228 = grantIsUncached ? release_ack_wait : _GEN_219;
  wire  _GEN_232 = grantIsCached & d_last;
  wire  _GEN_241 = grantIsCached ? release_ack_wait : _GEN_228;
  wire  _GEN_254 = _T_292 ? _GEN_241 : release_ack_wait;
  wire  tl_out__e_valid = grantIsRefill & ~dataArb_io_in_1_ready ? 1'h0 : auto_out_d_valid & d_first & grantIsCached &
    canAcceptCachedGrant;
  wire  _T_304 = auto_out_e_ready & tl_out__e_valid;
  wire [31:0] _dataArb_io_in_1_bits_addr_T_1 = {s2_vaddr[31:6], 6'h0};
  wire [31:0] _GEN_452 = {{20'd0}, d_address_inc};
  wire [31:0] _dataArb_io_in_1_bits_addr_T_2 = _dataArb_io_in_1_bits_addr_T_1 | _GEN_452;
  wire [3:0] _metaArb_io_in_3_bits_data_T_1 = {s2_write,_c_cat_T_49,auto_out_d_bits_param};
  wire [1:0] _metaArb_io_in_3_bits_data_T_11 = 4'h1 == _metaArb_io_in_3_bits_data_T_1 ? 2'h1 : 2'h0;
  wire [1:0] _metaArb_io_in_3_bits_data_T_13 = 4'h0 == _metaArb_io_in_3_bits_data_T_1 ? 2'h2 :
    _metaArb_io_in_3_bits_data_T_11;
  wire [1:0] _metaArb_io_in_3_bits_data_T_15 = 4'h4 == _metaArb_io_in_3_bits_data_T_1 ? 2'h2 :
    _metaArb_io_in_3_bits_data_T_13;
  wire [1:0] metaArb_io_in_3_bits_data_meta_state = 4'hc == _metaArb_io_in_3_bits_data_T_1 ? 2'h3 :
    _metaArb_io_in_3_bits_data_T_15;
  wire  _GEN_257 = auto_out_d_valid ? 1'h0 : _GEN_37;
  wire  _GEN_258 = auto_out_d_valid | auto_out_d_valid & grantIsRefill & canAcceptCachedGrant;
  wire  _GEN_259 = auto_out_d_valid ? 1'h0 : 1'h1;
  wire [9:0] counter1_1 = counter_1 - 10'h1;
  wire [9:0] _count_T_1 = ~counter1_1;
  wire [9:0] c_count = beats1_1 & _count_T_1;
  reg  s1_release_data_valid;
  wire  releaseRejected = s2_release_data_valid & ~_T_318;
  wire [10:0] _releaseDataBeat_T = {1'h0,c_count};
  wire [1:0] _releaseDataBeat_T_1 = {1'h0,s2_release_data_valid};
  wire [1:0] _GEN_453 = {{1'd0}, s1_release_data_valid};
  wire [1:0] _releaseDataBeat_T_3 = _GEN_453 + _releaseDataBeat_T_1;
  wire [1:0] _releaseDataBeat_T_4 = releaseRejected ? 2'h0 : _releaseDataBeat_T_3;
  wire [10:0] _GEN_454 = {{9'd0}, _releaseDataBeat_T_4};
  wire [10:0] releaseDataBeat = _releaseDataBeat_T + _GEN_454;
  wire  discard_line = s2_valid_flush_line & s2_req_size[1] | s2_flush_valid_pre_tag_ecc & flushing_req_size[1];
  wire [3:0] _release_state_T_13 = s2_victim_dirty & ~discard_line ? 4'h1 : 4'h6;
  wire [25:0] _probe_bits_T_2 = {s2_victim_tag,s2_req_addr[11:6]};
  wire [31:0] res_2_address = {_probe_bits_T_2, 6'h0};
  wire [3:0] _GEN_267 = s2_want_victimize ? _release_state_T_13 : release_state;
  wire [3:0] _release_state_T_14 = releaseDone ? 4'h7 : 4'h3;
  wire [3:0] _release_state_T_15 = releaseDone ? 4'h0 : 4'h5;
  wire [2:0] _GEN_278 = _T_324 ? s2_report_param : 3'h5;
  wire [3:0] _GEN_284 = _T_324 ? _release_state_T_14 : _release_state_T_15;
  wire [3:0] _GEN_286 = s2_prb_ack_data ? 4'h2 : _GEN_284;
  wire [2:0] _GEN_289 = s2_prb_ack_data ? 3'h5 : _GEN_278;
  wire [3:0] _GEN_307 = s2_probe ? _GEN_286 : _GEN_267;
  wire [2:0] _GEN_310 = s2_probe ? _GEN_289 : 3'h5;
  wire [32:0] _metaArb_io_in_6_bits_addr_T_3 = {1'h0,probe_bits_address};
  wire [3:0] _GEN_317 = metaArb_io_in_6_ready ? 4'h0 : _GEN_307;
  wire [32:0] _GEN_321 = release_state == 4'h4 ? _metaArb_io_in_6_bits_addr_T_3 : 33'h0;
  wire [3:0] _GEN_322 = release_state == 4'h4 ? _GEN_317 : _GEN_307;
  wire  _GEN_323 = release_state == 4'h4 & metaArb_io_in_6_ready;
  wire [3:0] _GEN_324 = releaseDone ? 4'h0 : _GEN_322;
  wire [3:0] _GEN_326 = release_state == 4'h5 ? _GEN_324 : _GEN_322;
  wire [3:0] _GEN_327 = releaseDone ? 4'h7 : _GEN_326;
  wire [2:0] _GEN_330 = release_state == 4'h3 ? s2_report_param : _GEN_310;
  wire [3:0] _GEN_336 = release_state == 4'h3 ? _GEN_327 : _GEN_326;
  wire [3:0] _GEN_337 = releaseDone ? 4'h7 : _GEN_336;
  wire [2:0] _GEN_339 = release_state == 4'h2 ? s2_report_param : _GEN_330;
  wire [3:0] _GEN_345 = release_state == 4'h2 ? _GEN_337 : _GEN_336;
  wire  _GEN_354 = _T_318 & c_first | _GEN_254;
  wire [1:0] newCoh_state = _T_333 ? voluntaryNewCoh_state : probeNewCoh_state;
  wire [11:0] _dataArb_io_in_2_bits_addr_T_1 = {probe_bits_address[11:6], 6'h0};
  wire [5:0] _dataArb_io_in_2_bits_addr_T_3 = {releaseDataBeat[3:0], 2'h0};
  wire [11:0] _GEN_467 = {{6'd0}, _dataArb_io_in_2_bits_addr_T_3};
  wire  _metaArb_io_in_4_valid_T_1 = release_state == 4'h7;
  wire [19:0] metaArb_io_in_4_bits_data_meta_tag = probe_bits_address[31:12];
  wire  _T_337 = metaArb_io_in_4_ready & metaArb_io_in_4_valid;
  reg  io_cpu_s2_xcpt_REG;
  reg  doUncachedResp;
  wire [15:0] io_cpu_resp_bits_data_shifted = get_a_mask_bit ? s2_data_corrected[31:16] : s2_data_corrected[15:0];
  wire  _io_cpu_resp_bits_data_T_3 = s2_req_signed & io_cpu_resp_bits_data_shifted[15];
  wire [15:0] _io_cpu_resp_bits_data_T_5 = _io_cpu_resp_bits_data_T_3 ? 16'hffff : 16'h0;
  wire [15:0] _io_cpu_resp_bits_data_T_7 = s2_req_size == 2'h1 ? _io_cpu_resp_bits_data_T_5 : s2_data_corrected[31:16];
  wire [31:0] _io_cpu_resp_bits_data_T_8 = {_io_cpu_resp_bits_data_T_7,io_cpu_resp_bits_data_shifted};
  wire [7:0] io_cpu_resp_bits_data_shifted_1 = get_a_mask_bit_1 ? _io_cpu_resp_bits_data_T_8[15:8] :
    _io_cpu_resp_bits_data_T_8[7:0];
  wire [7:0] io_cpu_resp_bits_data_zeroed_1 = _s2_write_T_3 ? 8'h0 : io_cpu_resp_bits_data_shifted_1;
  wire  _io_cpu_resp_bits_data_T_12 = s2_req_signed & io_cpu_resp_bits_data_zeroed_1[7];
  wire [23:0] _io_cpu_resp_bits_data_T_14 = _io_cpu_resp_bits_data_T_12 ? 24'hffffff : 24'h0;
  wire [23:0] _io_cpu_resp_bits_data_T_16 = s2_req_size == 2'h0 | _s2_write_T_3 ? _io_cpu_resp_bits_data_T_14 :
    _io_cpu_resp_bits_data_T_8[31:8];
  wire [31:0] _io_cpu_resp_bits_data_T_17 = {_io_cpu_resp_bits_data_T_16,io_cpu_resp_bits_data_zeroed_1};
  wire [31:0] _GEN_468 = {{31'd0}, s2_sc_fail};
  reg  REG;
  wire  _GEN_372 = REG | resetting;
  wire [8:0] flushCounterNext = flushCounter + 8'h1;
  wire  flushDone = flushCounterNext[8:6] == 3'h4;
  wire  _T_345 = s2_valid_masked & s2_cmd_flush_all;
  wire  _s1_flush_valid_T = metaArb_io_in_5_ready & metaArb_io_in_5_valid;
  wire  _metaArb_io_in_5_valid_T = ~flushed;
  wire [11:0] _metaArb_io_in_5_bits_addr_T_1 = {metaArb_io_in_5_bits_idx, 6'h0};
  wire  _GEN_373 = _metaArb_io_in_5_valid_T & _tl_out_a_valid_T_7 & _s2_valid_cached_miss_T_3 | flushing;
  wire  _GEN_386 = _T_345 ? _GEN_373 : flushing;
  wire  _GEN_399 = _T_284 & _s2_valid_cached_miss_T ? 1'h0 : flushed;
  wire  _GEN_400 = flushDone | _GEN_399;
  wire [8:0] _GEN_401 = s2_flush_valid_pre_tag_ecc ? flushCounterNext : {{1'd0}, flushCounter};
  wire  _GEN_402 = s2_flush_valid_pre_tag_ecc ? _GEN_400 : _GEN_399;
  wire [8:0] _GEN_405 = flushing ? _GEN_401 : {{1'd0}, flushCounter};
  wire  _GEN_406 = flushing ? _GEN_402 : _GEN_399;
  wire [8:0] _GEN_409 = resetting ? flushCounterNext : _GEN_405;
  reg [9:0] io_cpu_perf_release_counter;
  wire [9:0] io_cpu_perf_release_counter1 = io_cpu_perf_release_counter - 10'h1;
  wire  io_cpu_perf_release_first = io_cpu_perf_release_counter == 10'h0;
  wire  io_cpu_perf_release_last = io_cpu_perf_release_counter == 10'h1 | beats1_1 == 10'h0;
  wire  _T_369 = ~grantIsCached;
  wire  _GEN_481 = _T_292 & _T_369;
  OptimizationBarrier tlb_mpu_ppn_barrier (
    .io_x_ppn(tlb_mpu_ppn_barrier_io_x_ppn),
    .io_x_u(tlb_mpu_ppn_barrier_io_x_u),
    .io_x_ae_ptw(tlb_mpu_ppn_barrier_io_x_ae_ptw),
    .io_x_ae_final(tlb_mpu_ppn_barrier_io_x_ae_final),
    .io_x_pf(tlb_mpu_ppn_barrier_io_x_pf),
    .io_x_gf(tlb_mpu_ppn_barrier_io_x_gf),
    .io_x_sw(tlb_mpu_ppn_barrier_io_x_sw),
    .io_x_sx(tlb_mpu_ppn_barrier_io_x_sx),
    .io_x_sr(tlb_mpu_ppn_barrier_io_x_sr),
    .io_x_pw(tlb_mpu_ppn_barrier_io_x_pw),
    .io_x_px(tlb_mpu_ppn_barrier_io_x_px),
    .io_x_pr(tlb_mpu_ppn_barrier_io_x_pr),
    .io_x_ppp(tlb_mpu_ppn_barrier_io_x_ppp),
    .io_x_pal(tlb_mpu_ppn_barrier_io_x_pal),
    .io_x_paa(tlb_mpu_ppn_barrier_io_x_paa),
    .io_x_eff(tlb_mpu_ppn_barrier_io_x_eff),
    .io_x_c(tlb_mpu_ppn_barrier_io_x_c),
    .io_y_ppn(tlb_mpu_ppn_barrier_io_y_ppn),
    .io_y_u(tlb_mpu_ppn_barrier_io_y_u),
    .io_y_ae_ptw(tlb_mpu_ppn_barrier_io_y_ae_ptw),
    .io_y_ae_final(tlb_mpu_ppn_barrier_io_y_ae_final),
    .io_y_pf(tlb_mpu_ppn_barrier_io_y_pf),
    .io_y_gf(tlb_mpu_ppn_barrier_io_y_gf),
    .io_y_sw(tlb_mpu_ppn_barrier_io_y_sw),
    .io_y_sx(tlb_mpu_ppn_barrier_io_y_sx),
    .io_y_sr(tlb_mpu_ppn_barrier_io_y_sr),
    .io_y_pw(tlb_mpu_ppn_barrier_io_y_pw),
    .io_y_px(tlb_mpu_ppn_barrier_io_y_px),
    .io_y_pr(tlb_mpu_ppn_barrier_io_y_pr),
    .io_y_ppp(tlb_mpu_ppn_barrier_io_y_ppp),
    .io_y_pal(tlb_mpu_ppn_barrier_io_y_pal),
    .io_y_paa(tlb_mpu_ppn_barrier_io_y_paa),
    .io_y_eff(tlb_mpu_ppn_barrier_io_y_eff),
    .io_y_c(tlb_mpu_ppn_barrier_io_y_c)
  );
  PMPChecker tlb_pmp (
    .io_prv(tlb_pmp_io_prv),
    .io_pmp_0_cfg_l(tlb_pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(tlb_pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(tlb_pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(tlb_pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(tlb_pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(tlb_pmp_io_pmp_0_addr),
    .io_pmp_0_mask(tlb_pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(tlb_pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(tlb_pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(tlb_pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(tlb_pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(tlb_pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(tlb_pmp_io_pmp_1_addr),
    .io_pmp_1_mask(tlb_pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(tlb_pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(tlb_pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(tlb_pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(tlb_pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(tlb_pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(tlb_pmp_io_pmp_2_addr),
    .io_pmp_2_mask(tlb_pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(tlb_pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(tlb_pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(tlb_pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(tlb_pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(tlb_pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(tlb_pmp_io_pmp_3_addr),
    .io_pmp_3_mask(tlb_pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(tlb_pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(tlb_pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(tlb_pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(tlb_pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(tlb_pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(tlb_pmp_io_pmp_4_addr),
    .io_pmp_4_mask(tlb_pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(tlb_pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(tlb_pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(tlb_pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(tlb_pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(tlb_pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(tlb_pmp_io_pmp_5_addr),
    .io_pmp_5_mask(tlb_pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(tlb_pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(tlb_pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(tlb_pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(tlb_pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(tlb_pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(tlb_pmp_io_pmp_6_addr),
    .io_pmp_6_mask(tlb_pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(tlb_pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(tlb_pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(tlb_pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(tlb_pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(tlb_pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(tlb_pmp_io_pmp_7_addr),
    .io_pmp_7_mask(tlb_pmp_io_pmp_7_mask),
    .io_addr(tlb_pmp_io_addr),
    .io_r(tlb_pmp_io_r),
    .io_w(tlb_pmp_io_w),
    .io_x(tlb_pmp_io_x)
  );
  OptimizationBarrier tlb_entries_barrier (
    .io_x_ppn(tlb_entries_barrier_io_x_ppn),
    .io_x_u(tlb_entries_barrier_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_io_x_pf),
    .io_x_gf(tlb_entries_barrier_io_x_gf),
    .io_x_sw(tlb_entries_barrier_io_x_sw),
    .io_x_sx(tlb_entries_barrier_io_x_sx),
    .io_x_sr(tlb_entries_barrier_io_x_sr),
    .io_x_pw(tlb_entries_barrier_io_x_pw),
    .io_x_px(tlb_entries_barrier_io_x_px),
    .io_x_pr(tlb_entries_barrier_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_io_x_pal),
    .io_x_paa(tlb_entries_barrier_io_x_paa),
    .io_x_eff(tlb_entries_barrier_io_x_eff),
    .io_x_c(tlb_entries_barrier_io_x_c),
    .io_y_ppn(tlb_entries_barrier_io_y_ppn),
    .io_y_u(tlb_entries_barrier_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_io_y_pf),
    .io_y_gf(tlb_entries_barrier_io_y_gf),
    .io_y_sw(tlb_entries_barrier_io_y_sw),
    .io_y_sx(tlb_entries_barrier_io_y_sx),
    .io_y_sr(tlb_entries_barrier_io_y_sr),
    .io_y_pw(tlb_entries_barrier_io_y_pw),
    .io_y_px(tlb_entries_barrier_io_y_px),
    .io_y_pr(tlb_entries_barrier_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_io_y_pal),
    .io_y_paa(tlb_entries_barrier_io_y_paa),
    .io_y_eff(tlb_entries_barrier_io_y_eff),
    .io_y_c(tlb_entries_barrier_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_1 (
    .io_x_ppn(tlb_entries_barrier_1_io_x_ppn),
    .io_x_u(tlb_entries_barrier_1_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_1_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_1_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_1_io_x_pf),
    .io_x_gf(tlb_entries_barrier_1_io_x_gf),
    .io_x_sw(tlb_entries_barrier_1_io_x_sw),
    .io_x_sx(tlb_entries_barrier_1_io_x_sx),
    .io_x_sr(tlb_entries_barrier_1_io_x_sr),
    .io_x_pw(tlb_entries_barrier_1_io_x_pw),
    .io_x_px(tlb_entries_barrier_1_io_x_px),
    .io_x_pr(tlb_entries_barrier_1_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_1_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_1_io_x_pal),
    .io_x_paa(tlb_entries_barrier_1_io_x_paa),
    .io_x_eff(tlb_entries_barrier_1_io_x_eff),
    .io_x_c(tlb_entries_barrier_1_io_x_c),
    .io_y_ppn(tlb_entries_barrier_1_io_y_ppn),
    .io_y_u(tlb_entries_barrier_1_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_1_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_1_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_1_io_y_pf),
    .io_y_gf(tlb_entries_barrier_1_io_y_gf),
    .io_y_sw(tlb_entries_barrier_1_io_y_sw),
    .io_y_sx(tlb_entries_barrier_1_io_y_sx),
    .io_y_sr(tlb_entries_barrier_1_io_y_sr),
    .io_y_pw(tlb_entries_barrier_1_io_y_pw),
    .io_y_px(tlb_entries_barrier_1_io_y_px),
    .io_y_pr(tlb_entries_barrier_1_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_1_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_1_io_y_pal),
    .io_y_paa(tlb_entries_barrier_1_io_y_paa),
    .io_y_eff(tlb_entries_barrier_1_io_y_eff),
    .io_y_c(tlb_entries_barrier_1_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_2 (
    .io_x_ppn(tlb_entries_barrier_2_io_x_ppn),
    .io_x_u(tlb_entries_barrier_2_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_2_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_2_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_2_io_x_pf),
    .io_x_gf(tlb_entries_barrier_2_io_x_gf),
    .io_x_sw(tlb_entries_barrier_2_io_x_sw),
    .io_x_sx(tlb_entries_barrier_2_io_x_sx),
    .io_x_sr(tlb_entries_barrier_2_io_x_sr),
    .io_x_pw(tlb_entries_barrier_2_io_x_pw),
    .io_x_px(tlb_entries_barrier_2_io_x_px),
    .io_x_pr(tlb_entries_barrier_2_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_2_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_2_io_x_pal),
    .io_x_paa(tlb_entries_barrier_2_io_x_paa),
    .io_x_eff(tlb_entries_barrier_2_io_x_eff),
    .io_x_c(tlb_entries_barrier_2_io_x_c),
    .io_y_ppn(tlb_entries_barrier_2_io_y_ppn),
    .io_y_u(tlb_entries_barrier_2_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_2_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_2_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_2_io_y_pf),
    .io_y_gf(tlb_entries_barrier_2_io_y_gf),
    .io_y_sw(tlb_entries_barrier_2_io_y_sw),
    .io_y_sx(tlb_entries_barrier_2_io_y_sx),
    .io_y_sr(tlb_entries_barrier_2_io_y_sr),
    .io_y_pw(tlb_entries_barrier_2_io_y_pw),
    .io_y_px(tlb_entries_barrier_2_io_y_px),
    .io_y_pr(tlb_entries_barrier_2_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_2_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_2_io_y_pal),
    .io_y_paa(tlb_entries_barrier_2_io_y_paa),
    .io_y_eff(tlb_entries_barrier_2_io_y_eff),
    .io_y_c(tlb_entries_barrier_2_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_3 (
    .io_x_ppn(tlb_entries_barrier_3_io_x_ppn),
    .io_x_u(tlb_entries_barrier_3_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_3_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_3_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_3_io_x_pf),
    .io_x_gf(tlb_entries_barrier_3_io_x_gf),
    .io_x_sw(tlb_entries_barrier_3_io_x_sw),
    .io_x_sx(tlb_entries_barrier_3_io_x_sx),
    .io_x_sr(tlb_entries_barrier_3_io_x_sr),
    .io_x_pw(tlb_entries_barrier_3_io_x_pw),
    .io_x_px(tlb_entries_barrier_3_io_x_px),
    .io_x_pr(tlb_entries_barrier_3_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_3_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_3_io_x_pal),
    .io_x_paa(tlb_entries_barrier_3_io_x_paa),
    .io_x_eff(tlb_entries_barrier_3_io_x_eff),
    .io_x_c(tlb_entries_barrier_3_io_x_c),
    .io_y_ppn(tlb_entries_barrier_3_io_y_ppn),
    .io_y_u(tlb_entries_barrier_3_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_3_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_3_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_3_io_y_pf),
    .io_y_gf(tlb_entries_barrier_3_io_y_gf),
    .io_y_sw(tlb_entries_barrier_3_io_y_sw),
    .io_y_sx(tlb_entries_barrier_3_io_y_sx),
    .io_y_sr(tlb_entries_barrier_3_io_y_sr),
    .io_y_pw(tlb_entries_barrier_3_io_y_pw),
    .io_y_px(tlb_entries_barrier_3_io_y_px),
    .io_y_pr(tlb_entries_barrier_3_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_3_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_3_io_y_pal),
    .io_y_paa(tlb_entries_barrier_3_io_y_paa),
    .io_y_eff(tlb_entries_barrier_3_io_y_eff),
    .io_y_c(tlb_entries_barrier_3_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_4 (
    .io_x_ppn(tlb_entries_barrier_4_io_x_ppn),
    .io_x_u(tlb_entries_barrier_4_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_4_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_4_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_4_io_x_pf),
    .io_x_gf(tlb_entries_barrier_4_io_x_gf),
    .io_x_sw(tlb_entries_barrier_4_io_x_sw),
    .io_x_sx(tlb_entries_barrier_4_io_x_sx),
    .io_x_sr(tlb_entries_barrier_4_io_x_sr),
    .io_x_pw(tlb_entries_barrier_4_io_x_pw),
    .io_x_px(tlb_entries_barrier_4_io_x_px),
    .io_x_pr(tlb_entries_barrier_4_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_4_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_4_io_x_pal),
    .io_x_paa(tlb_entries_barrier_4_io_x_paa),
    .io_x_eff(tlb_entries_barrier_4_io_x_eff),
    .io_x_c(tlb_entries_barrier_4_io_x_c),
    .io_y_ppn(tlb_entries_barrier_4_io_y_ppn),
    .io_y_u(tlb_entries_barrier_4_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_4_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_4_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_4_io_y_pf),
    .io_y_gf(tlb_entries_barrier_4_io_y_gf),
    .io_y_sw(tlb_entries_barrier_4_io_y_sw),
    .io_y_sx(tlb_entries_barrier_4_io_y_sx),
    .io_y_sr(tlb_entries_barrier_4_io_y_sr),
    .io_y_pw(tlb_entries_barrier_4_io_y_pw),
    .io_y_px(tlb_entries_barrier_4_io_y_px),
    .io_y_pr(tlb_entries_barrier_4_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_4_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_4_io_y_pal),
    .io_y_paa(tlb_entries_barrier_4_io_y_paa),
    .io_y_eff(tlb_entries_barrier_4_io_y_eff),
    .io_y_c(tlb_entries_barrier_4_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_5 (
    .io_x_ppn(tlb_entries_barrier_5_io_x_ppn),
    .io_x_u(tlb_entries_barrier_5_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_5_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_5_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_5_io_x_pf),
    .io_x_gf(tlb_entries_barrier_5_io_x_gf),
    .io_x_sw(tlb_entries_barrier_5_io_x_sw),
    .io_x_sx(tlb_entries_barrier_5_io_x_sx),
    .io_x_sr(tlb_entries_barrier_5_io_x_sr),
    .io_x_pw(tlb_entries_barrier_5_io_x_pw),
    .io_x_px(tlb_entries_barrier_5_io_x_px),
    .io_x_pr(tlb_entries_barrier_5_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_5_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_5_io_x_pal),
    .io_x_paa(tlb_entries_barrier_5_io_x_paa),
    .io_x_eff(tlb_entries_barrier_5_io_x_eff),
    .io_x_c(tlb_entries_barrier_5_io_x_c),
    .io_y_ppn(tlb_entries_barrier_5_io_y_ppn),
    .io_y_u(tlb_entries_barrier_5_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_5_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_5_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_5_io_y_pf),
    .io_y_gf(tlb_entries_barrier_5_io_y_gf),
    .io_y_sw(tlb_entries_barrier_5_io_y_sw),
    .io_y_sx(tlb_entries_barrier_5_io_y_sx),
    .io_y_sr(tlb_entries_barrier_5_io_y_sr),
    .io_y_pw(tlb_entries_barrier_5_io_y_pw),
    .io_y_px(tlb_entries_barrier_5_io_y_px),
    .io_y_pr(tlb_entries_barrier_5_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_5_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_5_io_y_pal),
    .io_y_paa(tlb_entries_barrier_5_io_y_paa),
    .io_y_eff(tlb_entries_barrier_5_io_y_eff),
    .io_y_c(tlb_entries_barrier_5_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_6 (
    .io_x_ppn(tlb_entries_barrier_6_io_x_ppn),
    .io_x_u(tlb_entries_barrier_6_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_6_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_6_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_6_io_x_pf),
    .io_x_gf(tlb_entries_barrier_6_io_x_gf),
    .io_x_sw(tlb_entries_barrier_6_io_x_sw),
    .io_x_sx(tlb_entries_barrier_6_io_x_sx),
    .io_x_sr(tlb_entries_barrier_6_io_x_sr),
    .io_x_pw(tlb_entries_barrier_6_io_x_pw),
    .io_x_px(tlb_entries_barrier_6_io_x_px),
    .io_x_pr(tlb_entries_barrier_6_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_6_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_6_io_x_pal),
    .io_x_paa(tlb_entries_barrier_6_io_x_paa),
    .io_x_eff(tlb_entries_barrier_6_io_x_eff),
    .io_x_c(tlb_entries_barrier_6_io_x_c),
    .io_y_ppn(tlb_entries_barrier_6_io_y_ppn),
    .io_y_u(tlb_entries_barrier_6_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_6_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_6_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_6_io_y_pf),
    .io_y_gf(tlb_entries_barrier_6_io_y_gf),
    .io_y_sw(tlb_entries_barrier_6_io_y_sw),
    .io_y_sx(tlb_entries_barrier_6_io_y_sx),
    .io_y_sr(tlb_entries_barrier_6_io_y_sr),
    .io_y_pw(tlb_entries_barrier_6_io_y_pw),
    .io_y_px(tlb_entries_barrier_6_io_y_px),
    .io_y_pr(tlb_entries_barrier_6_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_6_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_6_io_y_pal),
    .io_y_paa(tlb_entries_barrier_6_io_y_paa),
    .io_y_eff(tlb_entries_barrier_6_io_y_eff),
    .io_y_c(tlb_entries_barrier_6_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_7 (
    .io_x_ppn(tlb_entries_barrier_7_io_x_ppn),
    .io_x_u(tlb_entries_barrier_7_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_7_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_7_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_7_io_x_pf),
    .io_x_gf(tlb_entries_barrier_7_io_x_gf),
    .io_x_sw(tlb_entries_barrier_7_io_x_sw),
    .io_x_sx(tlb_entries_barrier_7_io_x_sx),
    .io_x_sr(tlb_entries_barrier_7_io_x_sr),
    .io_x_pw(tlb_entries_barrier_7_io_x_pw),
    .io_x_px(tlb_entries_barrier_7_io_x_px),
    .io_x_pr(tlb_entries_barrier_7_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_7_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_7_io_x_pal),
    .io_x_paa(tlb_entries_barrier_7_io_x_paa),
    .io_x_eff(tlb_entries_barrier_7_io_x_eff),
    .io_x_c(tlb_entries_barrier_7_io_x_c),
    .io_y_ppn(tlb_entries_barrier_7_io_y_ppn),
    .io_y_u(tlb_entries_barrier_7_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_7_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_7_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_7_io_y_pf),
    .io_y_gf(tlb_entries_barrier_7_io_y_gf),
    .io_y_sw(tlb_entries_barrier_7_io_y_sw),
    .io_y_sx(tlb_entries_barrier_7_io_y_sx),
    .io_y_sr(tlb_entries_barrier_7_io_y_sr),
    .io_y_pw(tlb_entries_barrier_7_io_y_pw),
    .io_y_px(tlb_entries_barrier_7_io_y_px),
    .io_y_pr(tlb_entries_barrier_7_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_7_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_7_io_y_pal),
    .io_y_paa(tlb_entries_barrier_7_io_y_paa),
    .io_y_eff(tlb_entries_barrier_7_io_y_eff),
    .io_y_c(tlb_entries_barrier_7_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_8 (
    .io_x_ppn(tlb_entries_barrier_8_io_x_ppn),
    .io_x_u(tlb_entries_barrier_8_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_8_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_8_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_8_io_x_pf),
    .io_x_gf(tlb_entries_barrier_8_io_x_gf),
    .io_x_sw(tlb_entries_barrier_8_io_x_sw),
    .io_x_sx(tlb_entries_barrier_8_io_x_sx),
    .io_x_sr(tlb_entries_barrier_8_io_x_sr),
    .io_x_pw(tlb_entries_barrier_8_io_x_pw),
    .io_x_px(tlb_entries_barrier_8_io_x_px),
    .io_x_pr(tlb_entries_barrier_8_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_8_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_8_io_x_pal),
    .io_x_paa(tlb_entries_barrier_8_io_x_paa),
    .io_x_eff(tlb_entries_barrier_8_io_x_eff),
    .io_x_c(tlb_entries_barrier_8_io_x_c),
    .io_y_ppn(tlb_entries_barrier_8_io_y_ppn),
    .io_y_u(tlb_entries_barrier_8_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_8_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_8_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_8_io_y_pf),
    .io_y_gf(tlb_entries_barrier_8_io_y_gf),
    .io_y_sw(tlb_entries_barrier_8_io_y_sw),
    .io_y_sx(tlb_entries_barrier_8_io_y_sx),
    .io_y_sr(tlb_entries_barrier_8_io_y_sr),
    .io_y_pw(tlb_entries_barrier_8_io_y_pw),
    .io_y_px(tlb_entries_barrier_8_io_y_px),
    .io_y_pr(tlb_entries_barrier_8_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_8_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_8_io_y_pal),
    .io_y_paa(tlb_entries_barrier_8_io_y_paa),
    .io_y_eff(tlb_entries_barrier_8_io_y_eff),
    .io_y_c(tlb_entries_barrier_8_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_9 (
    .io_x_ppn(tlb_entries_barrier_9_io_x_ppn),
    .io_x_u(tlb_entries_barrier_9_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_9_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_9_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_9_io_x_pf),
    .io_x_gf(tlb_entries_barrier_9_io_x_gf),
    .io_x_sw(tlb_entries_barrier_9_io_x_sw),
    .io_x_sx(tlb_entries_barrier_9_io_x_sx),
    .io_x_sr(tlb_entries_barrier_9_io_x_sr),
    .io_x_pw(tlb_entries_barrier_9_io_x_pw),
    .io_x_px(tlb_entries_barrier_9_io_x_px),
    .io_x_pr(tlb_entries_barrier_9_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_9_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_9_io_x_pal),
    .io_x_paa(tlb_entries_barrier_9_io_x_paa),
    .io_x_eff(tlb_entries_barrier_9_io_x_eff),
    .io_x_c(tlb_entries_barrier_9_io_x_c),
    .io_y_ppn(tlb_entries_barrier_9_io_y_ppn),
    .io_y_u(tlb_entries_barrier_9_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_9_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_9_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_9_io_y_pf),
    .io_y_gf(tlb_entries_barrier_9_io_y_gf),
    .io_y_sw(tlb_entries_barrier_9_io_y_sw),
    .io_y_sx(tlb_entries_barrier_9_io_y_sx),
    .io_y_sr(tlb_entries_barrier_9_io_y_sr),
    .io_y_pw(tlb_entries_barrier_9_io_y_pw),
    .io_y_px(tlb_entries_barrier_9_io_y_px),
    .io_y_pr(tlb_entries_barrier_9_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_9_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_9_io_y_pal),
    .io_y_paa(tlb_entries_barrier_9_io_y_paa),
    .io_y_eff(tlb_entries_barrier_9_io_y_eff),
    .io_y_c(tlb_entries_barrier_9_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_10 (
    .io_x_ppn(tlb_entries_barrier_10_io_x_ppn),
    .io_x_u(tlb_entries_barrier_10_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_10_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_10_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_10_io_x_pf),
    .io_x_gf(tlb_entries_barrier_10_io_x_gf),
    .io_x_sw(tlb_entries_barrier_10_io_x_sw),
    .io_x_sx(tlb_entries_barrier_10_io_x_sx),
    .io_x_sr(tlb_entries_barrier_10_io_x_sr),
    .io_x_pw(tlb_entries_barrier_10_io_x_pw),
    .io_x_px(tlb_entries_barrier_10_io_x_px),
    .io_x_pr(tlb_entries_barrier_10_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_10_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_10_io_x_pal),
    .io_x_paa(tlb_entries_barrier_10_io_x_paa),
    .io_x_eff(tlb_entries_barrier_10_io_x_eff),
    .io_x_c(tlb_entries_barrier_10_io_x_c),
    .io_y_ppn(tlb_entries_barrier_10_io_y_ppn),
    .io_y_u(tlb_entries_barrier_10_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_10_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_10_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_10_io_y_pf),
    .io_y_gf(tlb_entries_barrier_10_io_y_gf),
    .io_y_sw(tlb_entries_barrier_10_io_y_sw),
    .io_y_sx(tlb_entries_barrier_10_io_y_sx),
    .io_y_sr(tlb_entries_barrier_10_io_y_sr),
    .io_y_pw(tlb_entries_barrier_10_io_y_pw),
    .io_y_px(tlb_entries_barrier_10_io_y_px),
    .io_y_pr(tlb_entries_barrier_10_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_10_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_10_io_y_pal),
    .io_y_paa(tlb_entries_barrier_10_io_y_paa),
    .io_y_eff(tlb_entries_barrier_10_io_y_eff),
    .io_y_c(tlb_entries_barrier_10_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_11 (
    .io_x_ppn(tlb_entries_barrier_11_io_x_ppn),
    .io_x_u(tlb_entries_barrier_11_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_11_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_11_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_11_io_x_pf),
    .io_x_gf(tlb_entries_barrier_11_io_x_gf),
    .io_x_sw(tlb_entries_barrier_11_io_x_sw),
    .io_x_sx(tlb_entries_barrier_11_io_x_sx),
    .io_x_sr(tlb_entries_barrier_11_io_x_sr),
    .io_x_pw(tlb_entries_barrier_11_io_x_pw),
    .io_x_px(tlb_entries_barrier_11_io_x_px),
    .io_x_pr(tlb_entries_barrier_11_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_11_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_11_io_x_pal),
    .io_x_paa(tlb_entries_barrier_11_io_x_paa),
    .io_x_eff(tlb_entries_barrier_11_io_x_eff),
    .io_x_c(tlb_entries_barrier_11_io_x_c),
    .io_y_ppn(tlb_entries_barrier_11_io_y_ppn),
    .io_y_u(tlb_entries_barrier_11_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_11_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_11_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_11_io_y_pf),
    .io_y_gf(tlb_entries_barrier_11_io_y_gf),
    .io_y_sw(tlb_entries_barrier_11_io_y_sw),
    .io_y_sx(tlb_entries_barrier_11_io_y_sx),
    .io_y_sr(tlb_entries_barrier_11_io_y_sr),
    .io_y_pw(tlb_entries_barrier_11_io_y_pw),
    .io_y_px(tlb_entries_barrier_11_io_y_px),
    .io_y_pr(tlb_entries_barrier_11_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_11_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_11_io_y_pal),
    .io_y_paa(tlb_entries_barrier_11_io_y_paa),
    .io_y_eff(tlb_entries_barrier_11_io_y_eff),
    .io_y_c(tlb_entries_barrier_11_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_12 (
    .io_x_ppn(tlb_entries_barrier_12_io_x_ppn),
    .io_x_u(tlb_entries_barrier_12_io_x_u),
    .io_x_ae_ptw(tlb_entries_barrier_12_io_x_ae_ptw),
    .io_x_ae_final(tlb_entries_barrier_12_io_x_ae_final),
    .io_x_pf(tlb_entries_barrier_12_io_x_pf),
    .io_x_gf(tlb_entries_barrier_12_io_x_gf),
    .io_x_sw(tlb_entries_barrier_12_io_x_sw),
    .io_x_sx(tlb_entries_barrier_12_io_x_sx),
    .io_x_sr(tlb_entries_barrier_12_io_x_sr),
    .io_x_pw(tlb_entries_barrier_12_io_x_pw),
    .io_x_px(tlb_entries_barrier_12_io_x_px),
    .io_x_pr(tlb_entries_barrier_12_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_12_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_12_io_x_pal),
    .io_x_paa(tlb_entries_barrier_12_io_x_paa),
    .io_x_eff(tlb_entries_barrier_12_io_x_eff),
    .io_x_c(tlb_entries_barrier_12_io_x_c),
    .io_y_ppn(tlb_entries_barrier_12_io_y_ppn),
    .io_y_u(tlb_entries_barrier_12_io_y_u),
    .io_y_ae_ptw(tlb_entries_barrier_12_io_y_ae_ptw),
    .io_y_ae_final(tlb_entries_barrier_12_io_y_ae_final),
    .io_y_pf(tlb_entries_barrier_12_io_y_pf),
    .io_y_gf(tlb_entries_barrier_12_io_y_gf),
    .io_y_sw(tlb_entries_barrier_12_io_y_sw),
    .io_y_sx(tlb_entries_barrier_12_io_y_sx),
    .io_y_sr(tlb_entries_barrier_12_io_y_sr),
    .io_y_pw(tlb_entries_barrier_12_io_y_pw),
    .io_y_px(tlb_entries_barrier_12_io_y_px),
    .io_y_pr(tlb_entries_barrier_12_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_12_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_12_io_y_pal),
    .io_y_paa(tlb_entries_barrier_12_io_y_paa),
    .io_y_eff(tlb_entries_barrier_12_io_y_eff),
    .io_y_c(tlb_entries_barrier_12_io_y_c)
  );
  OptimizationBarrier pma_checker_mpu_ppn_barrier (
    .io_x_ppn(pma_checker_mpu_ppn_barrier_io_x_ppn),
    .io_x_u(pma_checker_mpu_ppn_barrier_io_x_u),
    .io_x_ae_ptw(pma_checker_mpu_ppn_barrier_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_mpu_ppn_barrier_io_x_ae_final),
    .io_x_pf(pma_checker_mpu_ppn_barrier_io_x_pf),
    .io_x_gf(pma_checker_mpu_ppn_barrier_io_x_gf),
    .io_x_sw(pma_checker_mpu_ppn_barrier_io_x_sw),
    .io_x_sx(pma_checker_mpu_ppn_barrier_io_x_sx),
    .io_x_sr(pma_checker_mpu_ppn_barrier_io_x_sr),
    .io_x_pw(pma_checker_mpu_ppn_barrier_io_x_pw),
    .io_x_px(pma_checker_mpu_ppn_barrier_io_x_px),
    .io_x_pr(pma_checker_mpu_ppn_barrier_io_x_pr),
    .io_x_ppp(pma_checker_mpu_ppn_barrier_io_x_ppp),
    .io_x_pal(pma_checker_mpu_ppn_barrier_io_x_pal),
    .io_x_paa(pma_checker_mpu_ppn_barrier_io_x_paa),
    .io_x_eff(pma_checker_mpu_ppn_barrier_io_x_eff),
    .io_x_c(pma_checker_mpu_ppn_barrier_io_x_c),
    .io_y_ppn(pma_checker_mpu_ppn_barrier_io_y_ppn),
    .io_y_u(pma_checker_mpu_ppn_barrier_io_y_u),
    .io_y_ae_ptw(pma_checker_mpu_ppn_barrier_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_mpu_ppn_barrier_io_y_ae_final),
    .io_y_pf(pma_checker_mpu_ppn_barrier_io_y_pf),
    .io_y_gf(pma_checker_mpu_ppn_barrier_io_y_gf),
    .io_y_sw(pma_checker_mpu_ppn_barrier_io_y_sw),
    .io_y_sx(pma_checker_mpu_ppn_barrier_io_y_sx),
    .io_y_sr(pma_checker_mpu_ppn_barrier_io_y_sr),
    .io_y_pw(pma_checker_mpu_ppn_barrier_io_y_pw),
    .io_y_px(pma_checker_mpu_ppn_barrier_io_y_px),
    .io_y_pr(pma_checker_mpu_ppn_barrier_io_y_pr),
    .io_y_ppp(pma_checker_mpu_ppn_barrier_io_y_ppp),
    .io_y_pal(pma_checker_mpu_ppn_barrier_io_y_pal),
    .io_y_paa(pma_checker_mpu_ppn_barrier_io_y_paa),
    .io_y_eff(pma_checker_mpu_ppn_barrier_io_y_eff),
    .io_y_c(pma_checker_mpu_ppn_barrier_io_y_c)
  );
  PMPChecker pma_checker_pmp (
    .io_prv(pma_checker_pmp_io_prv),
    .io_pmp_0_cfg_l(pma_checker_pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pma_checker_pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pma_checker_pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pma_checker_pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pma_checker_pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pma_checker_pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pma_checker_pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pma_checker_pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pma_checker_pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pma_checker_pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pma_checker_pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pma_checker_pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pma_checker_pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pma_checker_pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pma_checker_pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pma_checker_pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pma_checker_pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pma_checker_pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pma_checker_pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pma_checker_pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pma_checker_pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pma_checker_pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pma_checker_pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pma_checker_pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pma_checker_pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pma_checker_pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pma_checker_pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pma_checker_pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pma_checker_pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pma_checker_pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pma_checker_pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pma_checker_pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pma_checker_pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pma_checker_pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pma_checker_pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pma_checker_pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pma_checker_pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pma_checker_pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pma_checker_pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pma_checker_pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pma_checker_pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pma_checker_pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pma_checker_pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pma_checker_pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pma_checker_pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pma_checker_pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pma_checker_pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pma_checker_pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pma_checker_pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pma_checker_pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pma_checker_pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pma_checker_pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pma_checker_pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pma_checker_pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pma_checker_pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pma_checker_pmp_io_pmp_7_mask),
    .io_addr(pma_checker_pmp_io_addr),
    .io_r(pma_checker_pmp_io_r),
    .io_w(pma_checker_pmp_io_w),
    .io_x(pma_checker_pmp_io_x)
  );
  OptimizationBarrier pma_checker_entries_barrier (
    .io_x_ppn(pma_checker_entries_barrier_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_1 (
    .io_x_ppn(pma_checker_entries_barrier_1_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_1_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_1_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_1_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_1_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_1_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_1_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_1_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_1_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_1_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_1_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_1_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_1_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_1_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_1_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_1_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_1_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_1_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_1_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_1_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_1_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_1_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_1_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_1_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_1_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_1_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_1_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_1_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_1_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_1_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_1_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_1_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_1_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_1_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_2 (
    .io_x_ppn(pma_checker_entries_barrier_2_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_2_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_2_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_2_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_2_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_2_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_2_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_2_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_2_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_2_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_2_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_2_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_2_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_2_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_2_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_2_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_2_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_2_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_2_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_2_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_2_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_2_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_2_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_2_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_2_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_2_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_2_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_2_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_2_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_2_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_2_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_2_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_2_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_2_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_3 (
    .io_x_ppn(pma_checker_entries_barrier_3_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_3_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_3_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_3_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_3_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_3_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_3_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_3_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_3_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_3_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_3_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_3_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_3_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_3_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_3_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_3_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_3_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_3_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_3_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_3_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_3_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_3_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_3_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_3_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_3_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_3_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_3_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_3_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_3_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_3_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_3_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_3_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_3_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_3_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_4 (
    .io_x_ppn(pma_checker_entries_barrier_4_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_4_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_4_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_4_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_4_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_4_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_4_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_4_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_4_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_4_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_4_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_4_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_4_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_4_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_4_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_4_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_4_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_4_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_4_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_4_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_4_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_4_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_4_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_4_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_4_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_4_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_4_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_4_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_4_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_4_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_4_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_4_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_4_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_4_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_5 (
    .io_x_ppn(pma_checker_entries_barrier_5_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_5_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_5_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_5_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_5_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_5_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_5_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_5_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_5_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_5_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_5_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_5_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_5_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_5_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_5_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_5_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_5_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_5_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_5_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_5_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_5_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_5_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_5_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_5_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_5_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_5_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_5_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_5_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_5_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_5_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_5_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_5_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_5_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_5_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_6 (
    .io_x_ppn(pma_checker_entries_barrier_6_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_6_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_6_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_6_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_6_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_6_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_6_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_6_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_6_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_6_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_6_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_6_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_6_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_6_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_6_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_6_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_6_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_6_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_6_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_6_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_6_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_6_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_6_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_6_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_6_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_6_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_6_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_6_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_6_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_6_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_6_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_6_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_6_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_6_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_7 (
    .io_x_ppn(pma_checker_entries_barrier_7_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_7_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_7_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_7_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_7_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_7_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_7_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_7_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_7_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_7_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_7_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_7_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_7_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_7_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_7_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_7_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_7_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_7_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_7_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_7_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_7_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_7_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_7_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_7_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_7_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_7_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_7_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_7_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_7_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_7_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_7_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_7_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_7_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_7_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_8 (
    .io_x_ppn(pma_checker_entries_barrier_8_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_8_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_8_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_8_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_8_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_8_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_8_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_8_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_8_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_8_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_8_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_8_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_8_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_8_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_8_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_8_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_8_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_8_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_8_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_8_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_8_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_8_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_8_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_8_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_8_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_8_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_8_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_8_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_8_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_8_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_8_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_8_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_8_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_8_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_9 (
    .io_x_ppn(pma_checker_entries_barrier_9_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_9_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_9_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_9_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_9_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_9_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_9_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_9_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_9_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_9_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_9_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_9_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_9_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_9_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_9_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_9_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_9_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_9_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_9_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_9_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_9_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_9_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_9_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_9_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_9_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_9_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_9_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_9_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_9_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_9_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_9_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_9_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_9_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_9_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_10 (
    .io_x_ppn(pma_checker_entries_barrier_10_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_10_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_10_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_10_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_10_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_10_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_10_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_10_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_10_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_10_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_10_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_10_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_10_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_10_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_10_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_10_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_10_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_10_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_10_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_10_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_10_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_10_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_10_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_10_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_10_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_10_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_10_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_10_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_10_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_10_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_10_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_10_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_10_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_10_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_11 (
    .io_x_ppn(pma_checker_entries_barrier_11_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_11_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_11_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_11_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_11_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_11_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_11_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_11_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_11_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_11_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_11_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_11_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_11_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_11_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_11_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_11_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_11_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_11_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_11_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_11_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_11_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_11_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_11_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_11_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_11_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_11_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_11_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_11_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_11_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_11_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_11_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_11_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_11_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_11_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_12 (
    .io_x_ppn(pma_checker_entries_barrier_12_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_12_io_x_u),
    .io_x_ae_ptw(pma_checker_entries_barrier_12_io_x_ae_ptw),
    .io_x_ae_final(pma_checker_entries_barrier_12_io_x_ae_final),
    .io_x_pf(pma_checker_entries_barrier_12_io_x_pf),
    .io_x_gf(pma_checker_entries_barrier_12_io_x_gf),
    .io_x_sw(pma_checker_entries_barrier_12_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_12_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_12_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_12_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_12_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_12_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_12_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_12_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_12_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_12_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_12_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_12_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_12_io_y_u),
    .io_y_ae_ptw(pma_checker_entries_barrier_12_io_y_ae_ptw),
    .io_y_ae_final(pma_checker_entries_barrier_12_io_y_ae_final),
    .io_y_pf(pma_checker_entries_barrier_12_io_y_pf),
    .io_y_gf(pma_checker_entries_barrier_12_io_y_gf),
    .io_y_sw(pma_checker_entries_barrier_12_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_12_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_12_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_12_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_12_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_12_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_12_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_12_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_12_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_12_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_12_io_y_c)
  );
  MaxPeriodFibonacciLFSR lfsr_prng (
    .clock(lfsr_prng_clock),
    .reset(lfsr_prng_reset),
    .io_increment(lfsr_prng_io_increment),
    .io_out_0(lfsr_prng_io_out_0),
    .io_out_1(lfsr_prng_io_out_1),
    .io_out_2(lfsr_prng_io_out_2),
    .io_out_3(lfsr_prng_io_out_3),
    .io_out_4(lfsr_prng_io_out_4),
    .io_out_5(lfsr_prng_io_out_5),
    .io_out_6(lfsr_prng_io_out_6),
    .io_out_7(lfsr_prng_io_out_7),
    .io_out_8(lfsr_prng_io_out_8),
    .io_out_9(lfsr_prng_io_out_9),
    .io_out_10(lfsr_prng_io_out_10),
    .io_out_11(lfsr_prng_io_out_11),
    .io_out_12(lfsr_prng_io_out_12),
    .io_out_13(lfsr_prng_io_out_13),
    .io_out_14(lfsr_prng_io_out_14),
    .io_out_15(lfsr_prng_io_out_15)
  );
  tag_array tag_array (
    .RW0_addr(tag_array_RW0_addr),
    .RW0_en(tag_array_RW0_en),
    .RW0_clk(tag_array_RW0_clk),
    .RW0_wmode(tag_array_RW0_wmode),
    .RW0_wdata_0(tag_array_RW0_wdata_0),
    .RW0_wdata_1(tag_array_RW0_wdata_1),
    .RW0_wdata_2(tag_array_RW0_wdata_2),
    .RW0_wdata_3(tag_array_RW0_wdata_3),
    .RW0_rdata_0(tag_array_RW0_rdata_0),
    .RW0_rdata_1(tag_array_RW0_rdata_1),
    .RW0_rdata_2(tag_array_RW0_rdata_2),
    .RW0_rdata_3(tag_array_RW0_rdata_3),
    .RW0_wmask_0(tag_array_RW0_wmask_0),
    .RW0_wmask_1(tag_array_RW0_wmask_1),
    .RW0_wmask_2(tag_array_RW0_wmask_2),
    .RW0_wmask_3(tag_array_RW0_wmask_3)
  );
  DCacheDataArray data (
    .clock(data_clock),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3)
  );
  AMOALU amoalu (
    .io_mask(amoalu_io_mask),
    .io_cmd(amoalu_io_cmd),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out)
  );
  assign tlb_io_req_ready = tlb_state == 2'h0;
  assign tlb_io_resp_miss = tlb__io_resp_miss_T_1 | tlb_multipleHits;
  assign tlb_io_resp_paddr = {tlb__ppn_T_48,tlb__mpu_physaddr_T};
  assign tlb_io_resp_pf_ld = |tlb__io_resp_pf_ld_T_1;
  assign tlb_io_resp_pf_st = |tlb__io_resp_pf_st_T_1;
  assign tlb_io_resp_ae_ld = |tlb__io_resp_ae_ld_T;
  assign tlb_io_resp_ae_st = |tlb__io_resp_ae_st_T;
  assign tlb_io_resp_ma_ld = tlb_misaligned & tlb_cmd_read;
  assign tlb_io_resp_ma_st = tlb_misaligned & tlb_cmd_write;
  assign tlb_io_resp_cacheable = |tlb__io_resp_cacheable_T;
  assign tlb_io_ptw_req_valid = tlb_state == 2'h1;
  assign tlb_io_ptw_req_bits_bits_addr = tlb_r_refill_tag;
  assign tlb_io_ptw_req_bits_bits_need_gpa = tlb_r_need_gpa;
  assign tlb_mpu_ppn_barrier_io_x_ppn = tlb_special_entry_data_0[40:21];
  assign tlb_mpu_ppn_barrier_io_x_u = tlb_special_entry_data_0[20];
  assign tlb_mpu_ppn_barrier_io_x_ae_ptw = tlb_special_entry_data_0[18];
  assign tlb_mpu_ppn_barrier_io_x_ae_final = tlb_special_entry_data_0[17];
  assign tlb_mpu_ppn_barrier_io_x_pf = tlb_special_entry_data_0[16];
  assign tlb_mpu_ppn_barrier_io_x_gf = tlb_special_entry_data_0[15];
  assign tlb_mpu_ppn_barrier_io_x_sw = tlb_special_entry_data_0[14];
  assign tlb_mpu_ppn_barrier_io_x_sx = tlb_special_entry_data_0[13];
  assign tlb_mpu_ppn_barrier_io_x_sr = tlb_special_entry_data_0[12];
  assign tlb_mpu_ppn_barrier_io_x_pw = tlb_special_entry_data_0[8];
  assign tlb_mpu_ppn_barrier_io_x_px = tlb_special_entry_data_0[7];
  assign tlb_mpu_ppn_barrier_io_x_pr = tlb_special_entry_data_0[6];
  assign tlb_mpu_ppn_barrier_io_x_ppp = tlb_special_entry_data_0[5];
  assign tlb_mpu_ppn_barrier_io_x_pal = tlb_special_entry_data_0[4];
  assign tlb_mpu_ppn_barrier_io_x_paa = tlb_special_entry_data_0[3];
  assign tlb_mpu_ppn_barrier_io_x_eff = tlb_special_entry_data_0[2];
  assign tlb_mpu_ppn_barrier_io_x_c = tlb_special_entry_data_0[1];
  assign tlb_pmp_io_prv = tlb_mpu_priv[1:0];
  assign tlb_pmp_io_pmp_0_cfg_l = tlb_io_ptw_pmp_0_cfg_l;
  assign tlb_pmp_io_pmp_0_cfg_a = tlb_io_ptw_pmp_0_cfg_a;
  assign tlb_pmp_io_pmp_0_cfg_x = tlb_io_ptw_pmp_0_cfg_x;
  assign tlb_pmp_io_pmp_0_cfg_w = tlb_io_ptw_pmp_0_cfg_w;
  assign tlb_pmp_io_pmp_0_cfg_r = tlb_io_ptw_pmp_0_cfg_r;
  assign tlb_pmp_io_pmp_0_addr = tlb_io_ptw_pmp_0_addr;
  assign tlb_pmp_io_pmp_0_mask = tlb_io_ptw_pmp_0_mask;
  assign tlb_pmp_io_pmp_1_cfg_l = tlb_io_ptw_pmp_1_cfg_l;
  assign tlb_pmp_io_pmp_1_cfg_a = tlb_io_ptw_pmp_1_cfg_a;
  assign tlb_pmp_io_pmp_1_cfg_x = tlb_io_ptw_pmp_1_cfg_x;
  assign tlb_pmp_io_pmp_1_cfg_w = tlb_io_ptw_pmp_1_cfg_w;
  assign tlb_pmp_io_pmp_1_cfg_r = tlb_io_ptw_pmp_1_cfg_r;
  assign tlb_pmp_io_pmp_1_addr = tlb_io_ptw_pmp_1_addr;
  assign tlb_pmp_io_pmp_1_mask = tlb_io_ptw_pmp_1_mask;
  assign tlb_pmp_io_pmp_2_cfg_l = tlb_io_ptw_pmp_2_cfg_l;
  assign tlb_pmp_io_pmp_2_cfg_a = tlb_io_ptw_pmp_2_cfg_a;
  assign tlb_pmp_io_pmp_2_cfg_x = tlb_io_ptw_pmp_2_cfg_x;
  assign tlb_pmp_io_pmp_2_cfg_w = tlb_io_ptw_pmp_2_cfg_w;
  assign tlb_pmp_io_pmp_2_cfg_r = tlb_io_ptw_pmp_2_cfg_r;
  assign tlb_pmp_io_pmp_2_addr = tlb_io_ptw_pmp_2_addr;
  assign tlb_pmp_io_pmp_2_mask = tlb_io_ptw_pmp_2_mask;
  assign tlb_pmp_io_pmp_3_cfg_l = tlb_io_ptw_pmp_3_cfg_l;
  assign tlb_pmp_io_pmp_3_cfg_a = tlb_io_ptw_pmp_3_cfg_a;
  assign tlb_pmp_io_pmp_3_cfg_x = tlb_io_ptw_pmp_3_cfg_x;
  assign tlb_pmp_io_pmp_3_cfg_w = tlb_io_ptw_pmp_3_cfg_w;
  assign tlb_pmp_io_pmp_3_cfg_r = tlb_io_ptw_pmp_3_cfg_r;
  assign tlb_pmp_io_pmp_3_addr = tlb_io_ptw_pmp_3_addr;
  assign tlb_pmp_io_pmp_3_mask = tlb_io_ptw_pmp_3_mask;
  assign tlb_pmp_io_pmp_4_cfg_l = tlb_io_ptw_pmp_4_cfg_l;
  assign tlb_pmp_io_pmp_4_cfg_a = tlb_io_ptw_pmp_4_cfg_a;
  assign tlb_pmp_io_pmp_4_cfg_x = tlb_io_ptw_pmp_4_cfg_x;
  assign tlb_pmp_io_pmp_4_cfg_w = tlb_io_ptw_pmp_4_cfg_w;
  assign tlb_pmp_io_pmp_4_cfg_r = tlb_io_ptw_pmp_4_cfg_r;
  assign tlb_pmp_io_pmp_4_addr = tlb_io_ptw_pmp_4_addr;
  assign tlb_pmp_io_pmp_4_mask = tlb_io_ptw_pmp_4_mask;
  assign tlb_pmp_io_pmp_5_cfg_l = tlb_io_ptw_pmp_5_cfg_l;
  assign tlb_pmp_io_pmp_5_cfg_a = tlb_io_ptw_pmp_5_cfg_a;
  assign tlb_pmp_io_pmp_5_cfg_x = tlb_io_ptw_pmp_5_cfg_x;
  assign tlb_pmp_io_pmp_5_cfg_w = tlb_io_ptw_pmp_5_cfg_w;
  assign tlb_pmp_io_pmp_5_cfg_r = tlb_io_ptw_pmp_5_cfg_r;
  assign tlb_pmp_io_pmp_5_addr = tlb_io_ptw_pmp_5_addr;
  assign tlb_pmp_io_pmp_5_mask = tlb_io_ptw_pmp_5_mask;
  assign tlb_pmp_io_pmp_6_cfg_l = tlb_io_ptw_pmp_6_cfg_l;
  assign tlb_pmp_io_pmp_6_cfg_a = tlb_io_ptw_pmp_6_cfg_a;
  assign tlb_pmp_io_pmp_6_cfg_x = tlb_io_ptw_pmp_6_cfg_x;
  assign tlb_pmp_io_pmp_6_cfg_w = tlb_io_ptw_pmp_6_cfg_w;
  assign tlb_pmp_io_pmp_6_cfg_r = tlb_io_ptw_pmp_6_cfg_r;
  assign tlb_pmp_io_pmp_6_addr = tlb_io_ptw_pmp_6_addr;
  assign tlb_pmp_io_pmp_6_mask = tlb_io_ptw_pmp_6_mask;
  assign tlb_pmp_io_pmp_7_cfg_l = tlb_io_ptw_pmp_7_cfg_l;
  assign tlb_pmp_io_pmp_7_cfg_a = tlb_io_ptw_pmp_7_cfg_a;
  assign tlb_pmp_io_pmp_7_cfg_x = tlb_io_ptw_pmp_7_cfg_x;
  assign tlb_pmp_io_pmp_7_cfg_w = tlb_io_ptw_pmp_7_cfg_w;
  assign tlb_pmp_io_pmp_7_cfg_r = tlb_io_ptw_pmp_7_cfg_r;
  assign tlb_pmp_io_pmp_7_addr = tlb_io_ptw_pmp_7_addr;
  assign tlb_pmp_io_pmp_7_mask = tlb_io_ptw_pmp_7_mask;
  assign tlb_pmp_io_addr = {tlb_mpu_ppn,tlb__mpu_physaddr_T};
  assign tlb_entries_barrier_io_x_ppn = tlb__GEN_609[40:21];
  assign tlb_entries_barrier_io_x_u = tlb__GEN_609[20];
  assign tlb_entries_barrier_io_x_ae_ptw = tlb__GEN_609[18];
  assign tlb_entries_barrier_io_x_ae_final = tlb__GEN_609[17];
  assign tlb_entries_barrier_io_x_pf = tlb__GEN_609[16];
  assign tlb_entries_barrier_io_x_gf = tlb__GEN_609[15];
  assign tlb_entries_barrier_io_x_sw = tlb__GEN_609[14];
  assign tlb_entries_barrier_io_x_sx = tlb__GEN_609[13];
  assign tlb_entries_barrier_io_x_sr = tlb__GEN_609[12];
  assign tlb_entries_barrier_io_x_pw = tlb__GEN_609[8];
  assign tlb_entries_barrier_io_x_px = tlb__GEN_609[7];
  assign tlb_entries_barrier_io_x_pr = tlb__GEN_609[6];
  assign tlb_entries_barrier_io_x_ppp = tlb__GEN_609[5];
  assign tlb_entries_barrier_io_x_pal = tlb__GEN_609[4];
  assign tlb_entries_barrier_io_x_paa = tlb__GEN_609[3];
  assign tlb_entries_barrier_io_x_eff = tlb__GEN_609[2];
  assign tlb_entries_barrier_io_x_c = tlb__GEN_609[1];
  assign tlb_entries_barrier_1_io_x_ppn = tlb__GEN_613[40:21];
  assign tlb_entries_barrier_1_io_x_u = tlb__GEN_613[20];
  assign tlb_entries_barrier_1_io_x_ae_ptw = tlb__GEN_613[18];
  assign tlb_entries_barrier_1_io_x_ae_final = tlb__GEN_613[17];
  assign tlb_entries_barrier_1_io_x_pf = tlb__GEN_613[16];
  assign tlb_entries_barrier_1_io_x_gf = tlb__GEN_613[15];
  assign tlb_entries_barrier_1_io_x_sw = tlb__GEN_613[14];
  assign tlb_entries_barrier_1_io_x_sx = tlb__GEN_613[13];
  assign tlb_entries_barrier_1_io_x_sr = tlb__GEN_613[12];
  assign tlb_entries_barrier_1_io_x_pw = tlb__GEN_613[8];
  assign tlb_entries_barrier_1_io_x_px = tlb__GEN_613[7];
  assign tlb_entries_barrier_1_io_x_pr = tlb__GEN_613[6];
  assign tlb_entries_barrier_1_io_x_ppp = tlb__GEN_613[5];
  assign tlb_entries_barrier_1_io_x_pal = tlb__GEN_613[4];
  assign tlb_entries_barrier_1_io_x_paa = tlb__GEN_613[3];
  assign tlb_entries_barrier_1_io_x_eff = tlb__GEN_613[2];
  assign tlb_entries_barrier_1_io_x_c = tlb__GEN_613[1];
  assign tlb_entries_barrier_2_io_x_ppn = tlb__GEN_617[40:21];
  assign tlb_entries_barrier_2_io_x_u = tlb__GEN_617[20];
  assign tlb_entries_barrier_2_io_x_ae_ptw = tlb__GEN_617[18];
  assign tlb_entries_barrier_2_io_x_ae_final = tlb__GEN_617[17];
  assign tlb_entries_barrier_2_io_x_pf = tlb__GEN_617[16];
  assign tlb_entries_barrier_2_io_x_gf = tlb__GEN_617[15];
  assign tlb_entries_barrier_2_io_x_sw = tlb__GEN_617[14];
  assign tlb_entries_barrier_2_io_x_sx = tlb__GEN_617[13];
  assign tlb_entries_barrier_2_io_x_sr = tlb__GEN_617[12];
  assign tlb_entries_barrier_2_io_x_pw = tlb__GEN_617[8];
  assign tlb_entries_barrier_2_io_x_px = tlb__GEN_617[7];
  assign tlb_entries_barrier_2_io_x_pr = tlb__GEN_617[6];
  assign tlb_entries_barrier_2_io_x_ppp = tlb__GEN_617[5];
  assign tlb_entries_barrier_2_io_x_pal = tlb__GEN_617[4];
  assign tlb_entries_barrier_2_io_x_paa = tlb__GEN_617[3];
  assign tlb_entries_barrier_2_io_x_eff = tlb__GEN_617[2];
  assign tlb_entries_barrier_2_io_x_c = tlb__GEN_617[1];
  assign tlb_entries_barrier_3_io_x_ppn = tlb__GEN_621[40:21];
  assign tlb_entries_barrier_3_io_x_u = tlb__GEN_621[20];
  assign tlb_entries_barrier_3_io_x_ae_ptw = tlb__GEN_621[18];
  assign tlb_entries_barrier_3_io_x_ae_final = tlb__GEN_621[17];
  assign tlb_entries_barrier_3_io_x_pf = tlb__GEN_621[16];
  assign tlb_entries_barrier_3_io_x_gf = tlb__GEN_621[15];
  assign tlb_entries_barrier_3_io_x_sw = tlb__GEN_621[14];
  assign tlb_entries_barrier_3_io_x_sx = tlb__GEN_621[13];
  assign tlb_entries_barrier_3_io_x_sr = tlb__GEN_621[12];
  assign tlb_entries_barrier_3_io_x_pw = tlb__GEN_621[8];
  assign tlb_entries_barrier_3_io_x_px = tlb__GEN_621[7];
  assign tlb_entries_barrier_3_io_x_pr = tlb__GEN_621[6];
  assign tlb_entries_barrier_3_io_x_ppp = tlb__GEN_621[5];
  assign tlb_entries_barrier_3_io_x_pal = tlb__GEN_621[4];
  assign tlb_entries_barrier_3_io_x_paa = tlb__GEN_621[3];
  assign tlb_entries_barrier_3_io_x_eff = tlb__GEN_621[2];
  assign tlb_entries_barrier_3_io_x_c = tlb__GEN_621[1];
  assign tlb_entries_barrier_4_io_x_ppn = tlb__GEN_625[40:21];
  assign tlb_entries_barrier_4_io_x_u = tlb__GEN_625[20];
  assign tlb_entries_barrier_4_io_x_ae_ptw = tlb__GEN_625[18];
  assign tlb_entries_barrier_4_io_x_ae_final = tlb__GEN_625[17];
  assign tlb_entries_barrier_4_io_x_pf = tlb__GEN_625[16];
  assign tlb_entries_barrier_4_io_x_gf = tlb__GEN_625[15];
  assign tlb_entries_barrier_4_io_x_sw = tlb__GEN_625[14];
  assign tlb_entries_barrier_4_io_x_sx = tlb__GEN_625[13];
  assign tlb_entries_barrier_4_io_x_sr = tlb__GEN_625[12];
  assign tlb_entries_barrier_4_io_x_pw = tlb__GEN_625[8];
  assign tlb_entries_barrier_4_io_x_px = tlb__GEN_625[7];
  assign tlb_entries_barrier_4_io_x_pr = tlb__GEN_625[6];
  assign tlb_entries_barrier_4_io_x_ppp = tlb__GEN_625[5];
  assign tlb_entries_barrier_4_io_x_pal = tlb__GEN_625[4];
  assign tlb_entries_barrier_4_io_x_paa = tlb__GEN_625[3];
  assign tlb_entries_barrier_4_io_x_eff = tlb__GEN_625[2];
  assign tlb_entries_barrier_4_io_x_c = tlb__GEN_625[1];
  assign tlb_entries_barrier_5_io_x_ppn = tlb__GEN_629[40:21];
  assign tlb_entries_barrier_5_io_x_u = tlb__GEN_629[20];
  assign tlb_entries_barrier_5_io_x_ae_ptw = tlb__GEN_629[18];
  assign tlb_entries_barrier_5_io_x_ae_final = tlb__GEN_629[17];
  assign tlb_entries_barrier_5_io_x_pf = tlb__GEN_629[16];
  assign tlb_entries_barrier_5_io_x_gf = tlb__GEN_629[15];
  assign tlb_entries_barrier_5_io_x_sw = tlb__GEN_629[14];
  assign tlb_entries_barrier_5_io_x_sx = tlb__GEN_629[13];
  assign tlb_entries_barrier_5_io_x_sr = tlb__GEN_629[12];
  assign tlb_entries_barrier_5_io_x_pw = tlb__GEN_629[8];
  assign tlb_entries_barrier_5_io_x_px = tlb__GEN_629[7];
  assign tlb_entries_barrier_5_io_x_pr = tlb__GEN_629[6];
  assign tlb_entries_barrier_5_io_x_ppp = tlb__GEN_629[5];
  assign tlb_entries_barrier_5_io_x_pal = tlb__GEN_629[4];
  assign tlb_entries_barrier_5_io_x_paa = tlb__GEN_629[3];
  assign tlb_entries_barrier_5_io_x_eff = tlb__GEN_629[2];
  assign tlb_entries_barrier_5_io_x_c = tlb__GEN_629[1];
  assign tlb_entries_barrier_6_io_x_ppn = tlb__GEN_633[40:21];
  assign tlb_entries_barrier_6_io_x_u = tlb__GEN_633[20];
  assign tlb_entries_barrier_6_io_x_ae_ptw = tlb__GEN_633[18];
  assign tlb_entries_barrier_6_io_x_ae_final = tlb__GEN_633[17];
  assign tlb_entries_barrier_6_io_x_pf = tlb__GEN_633[16];
  assign tlb_entries_barrier_6_io_x_gf = tlb__GEN_633[15];
  assign tlb_entries_barrier_6_io_x_sw = tlb__GEN_633[14];
  assign tlb_entries_barrier_6_io_x_sx = tlb__GEN_633[13];
  assign tlb_entries_barrier_6_io_x_sr = tlb__GEN_633[12];
  assign tlb_entries_barrier_6_io_x_pw = tlb__GEN_633[8];
  assign tlb_entries_barrier_6_io_x_px = tlb__GEN_633[7];
  assign tlb_entries_barrier_6_io_x_pr = tlb__GEN_633[6];
  assign tlb_entries_barrier_6_io_x_ppp = tlb__GEN_633[5];
  assign tlb_entries_barrier_6_io_x_pal = tlb__GEN_633[4];
  assign tlb_entries_barrier_6_io_x_paa = tlb__GEN_633[3];
  assign tlb_entries_barrier_6_io_x_eff = tlb__GEN_633[2];
  assign tlb_entries_barrier_6_io_x_c = tlb__GEN_633[1];
  assign tlb_entries_barrier_7_io_x_ppn = tlb__GEN_637[40:21];
  assign tlb_entries_barrier_7_io_x_u = tlb__GEN_637[20];
  assign tlb_entries_barrier_7_io_x_ae_ptw = tlb__GEN_637[18];
  assign tlb_entries_barrier_7_io_x_ae_final = tlb__GEN_637[17];
  assign tlb_entries_barrier_7_io_x_pf = tlb__GEN_637[16];
  assign tlb_entries_barrier_7_io_x_gf = tlb__GEN_637[15];
  assign tlb_entries_barrier_7_io_x_sw = tlb__GEN_637[14];
  assign tlb_entries_barrier_7_io_x_sx = tlb__GEN_637[13];
  assign tlb_entries_barrier_7_io_x_sr = tlb__GEN_637[12];
  assign tlb_entries_barrier_7_io_x_pw = tlb__GEN_637[8];
  assign tlb_entries_barrier_7_io_x_px = tlb__GEN_637[7];
  assign tlb_entries_barrier_7_io_x_pr = tlb__GEN_637[6];
  assign tlb_entries_barrier_7_io_x_ppp = tlb__GEN_637[5];
  assign tlb_entries_barrier_7_io_x_pal = tlb__GEN_637[4];
  assign tlb_entries_barrier_7_io_x_paa = tlb__GEN_637[3];
  assign tlb_entries_barrier_7_io_x_eff = tlb__GEN_637[2];
  assign tlb_entries_barrier_7_io_x_c = tlb__GEN_637[1];
  assign tlb_entries_barrier_8_io_x_ppn = tlb_superpage_entries_0_data_0[40:21];
  assign tlb_entries_barrier_8_io_x_u = tlb_superpage_entries_0_data_0[20];
  assign tlb_entries_barrier_8_io_x_ae_ptw = tlb_superpage_entries_0_data_0[18];
  assign tlb_entries_barrier_8_io_x_ae_final = tlb_superpage_entries_0_data_0[17];
  assign tlb_entries_barrier_8_io_x_pf = tlb_superpage_entries_0_data_0[16];
  assign tlb_entries_barrier_8_io_x_gf = tlb_superpage_entries_0_data_0[15];
  assign tlb_entries_barrier_8_io_x_sw = tlb_superpage_entries_0_data_0[14];
  assign tlb_entries_barrier_8_io_x_sx = tlb_superpage_entries_0_data_0[13];
  assign tlb_entries_barrier_8_io_x_sr = tlb_superpage_entries_0_data_0[12];
  assign tlb_entries_barrier_8_io_x_pw = tlb_superpage_entries_0_data_0[8];
  assign tlb_entries_barrier_8_io_x_px = tlb_superpage_entries_0_data_0[7];
  assign tlb_entries_barrier_8_io_x_pr = tlb_superpage_entries_0_data_0[6];
  assign tlb_entries_barrier_8_io_x_ppp = tlb_superpage_entries_0_data_0[5];
  assign tlb_entries_barrier_8_io_x_pal = tlb_superpage_entries_0_data_0[4];
  assign tlb_entries_barrier_8_io_x_paa = tlb_superpage_entries_0_data_0[3];
  assign tlb_entries_barrier_8_io_x_eff = tlb_superpage_entries_0_data_0[2];
  assign tlb_entries_barrier_8_io_x_c = tlb_superpage_entries_0_data_0[1];
  assign tlb_entries_barrier_9_io_x_ppn = tlb_superpage_entries_1_data_0[40:21];
  assign tlb_entries_barrier_9_io_x_u = tlb_superpage_entries_1_data_0[20];
  assign tlb_entries_barrier_9_io_x_ae_ptw = tlb_superpage_entries_1_data_0[18];
  assign tlb_entries_barrier_9_io_x_ae_final = tlb_superpage_entries_1_data_0[17];
  assign tlb_entries_barrier_9_io_x_pf = tlb_superpage_entries_1_data_0[16];
  assign tlb_entries_barrier_9_io_x_gf = tlb_superpage_entries_1_data_0[15];
  assign tlb_entries_barrier_9_io_x_sw = tlb_superpage_entries_1_data_0[14];
  assign tlb_entries_barrier_9_io_x_sx = tlb_superpage_entries_1_data_0[13];
  assign tlb_entries_barrier_9_io_x_sr = tlb_superpage_entries_1_data_0[12];
  assign tlb_entries_barrier_9_io_x_pw = tlb_superpage_entries_1_data_0[8];
  assign tlb_entries_barrier_9_io_x_px = tlb_superpage_entries_1_data_0[7];
  assign tlb_entries_barrier_9_io_x_pr = tlb_superpage_entries_1_data_0[6];
  assign tlb_entries_barrier_9_io_x_ppp = tlb_superpage_entries_1_data_0[5];
  assign tlb_entries_barrier_9_io_x_pal = tlb_superpage_entries_1_data_0[4];
  assign tlb_entries_barrier_9_io_x_paa = tlb_superpage_entries_1_data_0[3];
  assign tlb_entries_barrier_9_io_x_eff = tlb_superpage_entries_1_data_0[2];
  assign tlb_entries_barrier_9_io_x_c = tlb_superpage_entries_1_data_0[1];
  assign tlb_entries_barrier_10_io_x_ppn = tlb_superpage_entries_2_data_0[40:21];
  assign tlb_entries_barrier_10_io_x_u = tlb_superpage_entries_2_data_0[20];
  assign tlb_entries_barrier_10_io_x_ae_ptw = tlb_superpage_entries_2_data_0[18];
  assign tlb_entries_barrier_10_io_x_ae_final = tlb_superpage_entries_2_data_0[17];
  assign tlb_entries_barrier_10_io_x_pf = tlb_superpage_entries_2_data_0[16];
  assign tlb_entries_barrier_10_io_x_gf = tlb_superpage_entries_2_data_0[15];
  assign tlb_entries_barrier_10_io_x_sw = tlb_superpage_entries_2_data_0[14];
  assign tlb_entries_barrier_10_io_x_sx = tlb_superpage_entries_2_data_0[13];
  assign tlb_entries_barrier_10_io_x_sr = tlb_superpage_entries_2_data_0[12];
  assign tlb_entries_barrier_10_io_x_pw = tlb_superpage_entries_2_data_0[8];
  assign tlb_entries_barrier_10_io_x_px = tlb_superpage_entries_2_data_0[7];
  assign tlb_entries_barrier_10_io_x_pr = tlb_superpage_entries_2_data_0[6];
  assign tlb_entries_barrier_10_io_x_ppp = tlb_superpage_entries_2_data_0[5];
  assign tlb_entries_barrier_10_io_x_pal = tlb_superpage_entries_2_data_0[4];
  assign tlb_entries_barrier_10_io_x_paa = tlb_superpage_entries_2_data_0[3];
  assign tlb_entries_barrier_10_io_x_eff = tlb_superpage_entries_2_data_0[2];
  assign tlb_entries_barrier_10_io_x_c = tlb_superpage_entries_2_data_0[1];
  assign tlb_entries_barrier_11_io_x_ppn = tlb_superpage_entries_3_data_0[40:21];
  assign tlb_entries_barrier_11_io_x_u = tlb_superpage_entries_3_data_0[20];
  assign tlb_entries_barrier_11_io_x_ae_ptw = tlb_superpage_entries_3_data_0[18];
  assign tlb_entries_barrier_11_io_x_ae_final = tlb_superpage_entries_3_data_0[17];
  assign tlb_entries_barrier_11_io_x_pf = tlb_superpage_entries_3_data_0[16];
  assign tlb_entries_barrier_11_io_x_gf = tlb_superpage_entries_3_data_0[15];
  assign tlb_entries_barrier_11_io_x_sw = tlb_superpage_entries_3_data_0[14];
  assign tlb_entries_barrier_11_io_x_sx = tlb_superpage_entries_3_data_0[13];
  assign tlb_entries_barrier_11_io_x_sr = tlb_superpage_entries_3_data_0[12];
  assign tlb_entries_barrier_11_io_x_pw = tlb_superpage_entries_3_data_0[8];
  assign tlb_entries_barrier_11_io_x_px = tlb_superpage_entries_3_data_0[7];
  assign tlb_entries_barrier_11_io_x_pr = tlb_superpage_entries_3_data_0[6];
  assign tlb_entries_barrier_11_io_x_ppp = tlb_superpage_entries_3_data_0[5];
  assign tlb_entries_barrier_11_io_x_pal = tlb_superpage_entries_3_data_0[4];
  assign tlb_entries_barrier_11_io_x_paa = tlb_superpage_entries_3_data_0[3];
  assign tlb_entries_barrier_11_io_x_eff = tlb_superpage_entries_3_data_0[2];
  assign tlb_entries_barrier_11_io_x_c = tlb_superpage_entries_3_data_0[1];
  assign tlb_entries_barrier_12_io_x_ppn = tlb_special_entry_data_0[40:21];
  assign tlb_entries_barrier_12_io_x_u = tlb_special_entry_data_0[20];
  assign tlb_entries_barrier_12_io_x_ae_ptw = tlb_special_entry_data_0[18];
  assign tlb_entries_barrier_12_io_x_ae_final = tlb_special_entry_data_0[17];
  assign tlb_entries_barrier_12_io_x_pf = tlb_special_entry_data_0[16];
  assign tlb_entries_barrier_12_io_x_gf = tlb_special_entry_data_0[15];
  assign tlb_entries_barrier_12_io_x_sw = tlb_special_entry_data_0[14];
  assign tlb_entries_barrier_12_io_x_sx = tlb_special_entry_data_0[13];
  assign tlb_entries_barrier_12_io_x_sr = tlb_special_entry_data_0[12];
  assign tlb_entries_barrier_12_io_x_pw = tlb_special_entry_data_0[8];
  assign tlb_entries_barrier_12_io_x_px = tlb_special_entry_data_0[7];
  assign tlb_entries_barrier_12_io_x_pr = tlb_special_entry_data_0[6];
  assign tlb_entries_barrier_12_io_x_ppp = tlb_special_entry_data_0[5];
  assign tlb_entries_barrier_12_io_x_pal = tlb_special_entry_data_0[4];
  assign tlb_entries_barrier_12_io_x_paa = tlb_special_entry_data_0[3];
  assign tlb_entries_barrier_12_io_x_eff = tlb_special_entry_data_0[2];
  assign tlb_entries_barrier_12_io_x_c = tlb_special_entry_data_0[1];
  assign pma_checker_mpu_ppn_barrier_io_x_ppn = 20'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_u = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_ae_ptw = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_ae_final = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_pf = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_gf = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_sw = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_sx = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_sr = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_pw = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_px = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_pr = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_ppp = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_pal = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_paa = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_eff = 1'h0;
  assign pma_checker_mpu_ppn_barrier_io_x_c = 1'h0;
  assign pma_checker_pmp_io_prv = 2'h1;
  assign pma_checker_pmp_io_pmp_0_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_0_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_0_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_0_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_0_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_0_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_0_mask = 32'h0;
  assign pma_checker_pmp_io_pmp_1_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_1_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_1_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_1_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_1_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_1_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_1_mask = 32'h0;
  assign pma_checker_pmp_io_pmp_2_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_2_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_2_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_2_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_2_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_2_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_2_mask = 32'h0;
  assign pma_checker_pmp_io_pmp_3_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_3_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_3_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_3_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_3_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_3_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_3_mask = 32'h0;
  assign pma_checker_pmp_io_pmp_4_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_4_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_4_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_4_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_4_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_4_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_4_mask = 32'h0;
  assign pma_checker_pmp_io_pmp_5_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_5_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_5_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_5_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_5_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_5_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_5_mask = 32'h0;
  assign pma_checker_pmp_io_pmp_6_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_6_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_6_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_6_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_6_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_6_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_6_mask = 32'h0;
  assign pma_checker_pmp_io_pmp_7_cfg_l = 1'h0;
  assign pma_checker_pmp_io_pmp_7_cfg_a = 2'h0;
  assign pma_checker_pmp_io_pmp_7_cfg_x = 1'h0;
  assign pma_checker_pmp_io_pmp_7_cfg_w = 1'h0;
  assign pma_checker_pmp_io_pmp_7_cfg_r = 1'h0;
  assign pma_checker_pmp_io_pmp_7_addr = 30'h0;
  assign pma_checker_pmp_io_pmp_7_mask = 32'h0;
  assign pma_checker_pmp_io_addr = 32'h0;
  assign pma_checker_entries_barrier_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_1_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_1_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_2_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_2_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_3_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_3_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_4_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_4_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_5_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_5_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_6_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_6_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_7_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_7_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_8_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_8_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_9_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_9_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_10_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_10_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_11_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_11_io_x_c = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_ppn = 20'h0;
  assign pma_checker_entries_barrier_12_io_x_u = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_ae_ptw = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_ae_final = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_pf = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_gf = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_sw = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_sx = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_sr = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_pw = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_px = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_pr = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_ppp = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_pal = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_paa = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_eff = 1'h0;
  assign pma_checker_entries_barrier_12_io_x_c = 1'h0;
  assign metaArb_io_in_4_ready = ~metaArb__grant_T_2;
  assign metaArb_io_in_5_ready = ~metaArb__grant_T_3;
  assign metaArb_io_in_6_ready = ~metaArb__grant_T_4;
  assign metaArb_io_in_7_ready = ~metaArb__grant_T_5;
  assign metaArb_io_out_valid = metaArb__io_out_valid_T | metaArb_io_in_7_valid;
  assign metaArb_io_out_bits_write = metaArb_io_in_0_valid | metaArb__GEN_25;
  assign metaArb_io_out_bits_addr = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_addr : metaArb__GEN_26;
  assign metaArb_io_out_bits_idx = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_idx : metaArb__GEN_27;
  assign metaArb_io_out_bits_way_en = metaArb_io_in_0_valid ? 4'hf : metaArb__GEN_28;
  assign metaArb_io_out_bits_data = metaArb_io_in_0_valid ? 22'h0 : metaArb__GEN_29;
  assign dataArb_io_in_1_ready = ~dataArb_io_in_0_valid;
  assign dataArb_io_in_2_ready = ~dataArb__grant_T;
  assign dataArb_io_in_3_ready = ~dataArb__grant_T_1;
  assign dataArb_io_out_valid = dataArb__io_out_valid_T | dataArb_io_in_3_valid;
  assign dataArb_io_out_bits_addr = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_addr : dataArb__GEN_8;
  assign dataArb_io_out_bits_write = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_write : dataArb__GEN_9;
  assign dataArb_io_out_bits_wdata = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_wdata : dataArb__GEN_10;
  assign dataArb_io_out_bits_eccMask = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_eccMask : 4'hf;
  assign dataArb_io_out_bits_way_en = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_way_en : dataArb__GEN_13;
  assign auto_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12;
  assign auto_out_a_bits_opcode = _s2_valid_cached_miss_T ? 3'h6 : _tl_out_a_bits_T_8_opcode;
  assign auto_out_a_bits_param = _s2_valid_cached_miss_T ? tl_out_a_bits_a_param : _tl_out_a_bits_T_8_param;
  assign auto_out_a_bits_size = _s2_valid_cached_miss_T ? 4'h6 : _tl_out_a_bits_T_8_size;
  assign auto_out_a_bits_source = _s2_valid_cached_miss_T ? 1'h0 : _tl_out_a_bits_T_8_source;
  assign auto_out_a_bits_address = _s2_valid_cached_miss_T ? acquire_address : _tl_out_a_bits_T_8_address;
  assign auto_out_a_bits_mask = _s2_valid_cached_miss_T ? 4'hf : _tl_out_a_bits_T_8_mask;
  assign auto_out_a_bits_data = _s2_valid_cached_miss_T ? 32'h0 : _tl_out_a_bits_T_8_data;
  assign auto_out_c_valid = release_state == 4'h3 | _GEN_325;
  assign auto_out_c_bits_opcode = _T_333 ? _GEN_346 : _GEN_338;
  assign auto_out_c_bits_param = _T_333 ? s2_shrink_param : _GEN_339;
  assign auto_out_c_bits_size = _T_333 ? 4'h6 : 4'h0;
  assign auto_out_c_bits_address = probe_bits_address;
  assign auto_out_c_bits_data = {s2_data_corrected_hi,s2_data_corrected_lo};
  assign auto_out_d_ready = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? 1'h0 : _GEN_256;
  assign auto_out_e_valid = grantIsRefill & ~dataArb_io_in_1_ready ? 1'h0 : auto_out_d_valid & d_first & grantIsCached
     & canAcceptCachedGrant;
  assign auto_out_e_bits_sink = auto_out_d_bits_sink;
  assign io_cpu_req_ready = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? _GEN_257 : _GEN_37;
  assign io_cpu_s2_nack = s2_valid_no_xcpt & ~s2_dont_nack_uncached & ~s2_dont_nack_misc & ~
    s2_valid_hit_pre_data_ecc_and_waw;
  assign io_cpu_resp_valid = s2_valid_hit_pre_data_ecc_and_waw | doUncachedResp;
  assign io_cpu_resp_bits_addr = doUncachedResp ? s2_uncached_resp_addr : s2_req_addr;
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_cmd = s2_req_cmd;
  assign io_cpu_resp_bits_size = s2_req_size;
  assign io_cpu_resp_bits_signed = s2_req_signed;
  assign io_cpu_resp_bits_dprv = s2_req_dprv;
  assign io_cpu_resp_bits_dv = 1'h0;
  assign io_cpu_resp_bits_data = _io_cpu_resp_bits_data_T_17 | _GEN_468;
  assign io_cpu_resp_bits_mask = 4'h0;
  assign io_cpu_resp_bits_replay = doUncachedResp;
  assign io_cpu_resp_bits_has_data = _s2_read_T_6 | _s2_write_T_21;
  assign io_cpu_resp_bits_data_word_bypass = {s2_data_corrected_hi,s2_data_corrected_lo};
  assign io_cpu_resp_bits_data_raw = {s2_data_corrected_hi,s2_data_corrected_lo};
  assign io_cpu_resp_bits_store_data = pstore1_data;
  assign io_cpu_replay_next = _T_292 & grantIsUncachedData;
  assign io_cpu_s2_xcpt_ma_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_ld;
  assign io_cpu_s2_xcpt_ma_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_st;
  assign io_cpu_s2_xcpt_pf_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_ld;
  assign io_cpu_s2_xcpt_pf_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_st;
  assign io_cpu_s2_xcpt_gf_ld = 1'h0;
  assign io_cpu_s2_xcpt_gf_st = 1'h0;
  assign io_cpu_s2_xcpt_ae_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_ld;
  assign io_cpu_s2_xcpt_ae_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_st;
  assign io_cpu_ordered = ~(s1_valid | s2_valid | cached_grant_wait | _s2_valid_cached_miss_T_2);
  assign io_cpu_perf_release = io_cpu_perf_release_last & _T_318;
  assign io_cpu_perf_grant = auto_out_d_valid & d_last;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr;
  assign io_ptw_req_bits_bits_need_gpa = tlb_io_ptw_req_bits_bits_need_gpa;
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid_masked & s1_cmd_uses_tlb;
  assign tlb_io_req_bits_vaddr = s1_tlb_req_vaddr;
  assign tlb_io_req_bits_passthrough = s1_tlb_req_passthrough;
  assign tlb_io_req_bits_size = s1_tlb_req_size;
  assign tlb_io_req_bits_cmd = s1_tlb_req_cmd;
  assign tlb_io_req_bits_prv = s1_tlb_req_prv;
  assign tlb_io_sfence_valid = s1_valid_masked & s1_sfence;
  assign tlb_io_sfence_bits_rs1 = s1_req_size[0];
  assign tlb_io_sfence_bits_rs2 = s1_req_size[1];
  assign tlb_io_sfence_bits_addr = s1_req_addr;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_ae_ptw = io_ptw_resp_bits_ae_ptw;
  assign tlb_io_ptw_resp_bits_ae_final = io_ptw_resp_bits_ae_final;
  assign tlb_io_ptw_resp_bits_pf = io_ptw_resp_bits_pf;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a;
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g;
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u;
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x;
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level;
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous;
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_sum = io_ptw_status_sum;
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr;
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask;
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr;
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask;
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr;
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask;
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr;
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask;
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr;
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask;
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr;
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask;
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr;
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask;
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr;
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask;
  assign lfsr_prng_clock = clock;
  assign lfsr_prng_reset = reset;
  assign lfsr_prng_io_increment = _T_292 & _GEN_232;
  assign metaArb_io_in_0_valid = resetting;
  assign metaArb_io_in_0_bits_addr = metaArb_io_in_5_bits_addr;
  assign metaArb_io_in_0_bits_idx = metaArb_io_in_5_bits_idx;
  assign metaArb_io_in_2_valid = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta;
  assign metaArb_io_in_2_bits_addr = {io_cpu_req_bits_addr[31:12],s2_vaddr[11:0]};
  assign metaArb_io_in_2_bits_idx = s2_vaddr[11:6];
  assign metaArb_io_in_2_bits_way_en = s2_hit_valid ? s2_hit_way : s2_victim_way;
  assign metaArb_io_in_2_bits_data = {s2_grow_param,metaArb_io_in_2_bits_data_meta_tag};
  assign metaArb_io_in_3_valid = grantIsCached & d_done & ~auto_out_d_bits_denied;
  assign metaArb_io_in_3_bits_addr = {io_cpu_req_bits_addr[31:12],s2_vaddr[11:0]};
  assign metaArb_io_in_3_bits_idx = s2_vaddr[11:6];
  assign metaArb_io_in_3_bits_way_en = refill_way;
  assign metaArb_io_in_3_bits_data = {metaArb_io_in_3_bits_data_meta_state,metaArb_io_in_2_bits_data_meta_tag};
  assign metaArb_io_in_4_valid = _T_330 | _metaArb_io_in_4_valid_T_1;
  assign metaArb_io_in_4_bits_addr = {io_cpu_req_bits_addr[31:12],probe_bits_address[11:0]};
  assign metaArb_io_in_4_bits_idx = probe_bits_address[11:6];
  assign metaArb_io_in_4_bits_way_en = _T_333 ? s2_victim_or_hit_way : s2_probe_way;
  assign metaArb_io_in_4_bits_data = {newCoh_state,metaArb_io_in_4_bits_data_meta_tag};
  assign metaArb_io_in_5_valid = flushing & ~flushed;
  assign metaArb_io_in_5_bits_addr = {io_cpu_req_bits_addr[31:12],_metaArb_io_in_5_bits_addr_T_1};
  assign metaArb_io_in_5_bits_idx = flushCounter[5:0];
  assign metaArb_io_in_5_bits_way_en = metaArb_io_in_4_bits_way_en;
  assign metaArb_io_in_5_bits_data = metaArb_io_in_4_bits_data;
  assign metaArb_io_in_6_valid = release_state == 4'h4;
  assign metaArb_io_in_6_bits_addr = _GEN_321[31:0];
  assign metaArb_io_in_6_bits_idx = release_state == 4'h4 ? probe_bits_address[11:6] : 6'h0;
  assign metaArb_io_in_6_bits_way_en = metaArb_io_in_4_bits_way_en;
  assign metaArb_io_in_6_bits_data = metaArb_io_in_4_bits_data;
  assign metaArb_io_in_7_valid = io_cpu_req_valid;
  assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr;
  assign metaArb_io_in_7_bits_idx = dataArb_io_in_3_bits_addr[11:6];
  assign metaArb_io_in_7_bits_way_en = metaArb_io_in_4_bits_way_en;
  assign metaArb_io_in_7_bits_data = metaArb_io_in_4_bits_data;
  assign tag_array_RW0_clk = clock;
  assign tag_array_RW0_wdata_0 = metaArb_io_out_bits_data;
  assign tag_array_RW0_wdata_1 = metaArb_io_out_bits_data;
  assign tag_array_RW0_wdata_2 = metaArb_io_out_bits_data;
  assign tag_array_RW0_wdata_3 = metaArb_io_out_bits_data;
  assign tag_array_RW0_wmask_0 = metaArb_io_out_bits_way_en[0];
  assign tag_array_RW0_wmask_1 = metaArb_io_out_bits_way_en[1];
  assign tag_array_RW0_wmask_2 = metaArb_io_out_bits_way_en[2];
  assign tag_array_RW0_wmask_3 = metaArb_io_out_bits_way_en[3];
  assign data_clock = clock;
  assign data_io_req_valid = dataArb_io_out_valid;
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr;
  assign data_io_req_bits_write = dataArb_io_out_bits_write;
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata;
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask;
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en;
  assign dataArb_io_in_0_valid = pstore_drain_structural | _pstore_drain_T_10;
  assign dataArb_io_in_0_bits_addr = _dataArb_io_in_0_bits_addr_T[11:0];
  assign dataArb_io_in_0_bits_write = pstore_drain_structural | _pstore_drain_T_10;
  assign dataArb_io_in_0_bits_wdata = {dataArb_io_in_0_bits_wdata_hi,dataArb_io_in_0_bits_wdata_lo};
  assign dataArb_io_in_0_bits_eccMask = {dataArb_io_in_0_bits_eccMask_hi,dataArb_io_in_0_bits_eccMask_lo};
  assign dataArb_io_in_0_bits_way_en = pstore2_valid ? pstore2_way : pstore1_way;
  assign dataArb_io_in_1_valid = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? _GEN_258 : auto_out_d_valid &
    grantIsRefill & canAcceptCachedGrant;
  assign dataArb_io_in_1_bits_addr = _dataArb_io_in_1_bits_addr_T_2[11:0];
  assign dataArb_io_in_1_bits_write = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? _GEN_259 : 1'h1;
  assign dataArb_io_in_1_bits_wdata = {tl_d_data_encoded_hi,tl_d_data_encoded_lo};
  assign dataArb_io_in_1_bits_way_en = refill_way;
  assign dataArb_io_in_2_valid = inWriteback & releaseDataBeat < 11'h10;
  assign dataArb_io_in_2_bits_addr = _dataArb_io_in_2_bits_addr_T_1 | _GEN_467;
  assign dataArb_io_in_2_bits_wdata = dataArb_io_in_1_bits_wdata;
  assign dataArb_io_in_3_valid = io_cpu_req_valid & res;
  assign dataArb_io_in_3_bits_addr = _dataArb_io_in_3_bits_addr_T_2[11:0];
  assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata;
  assign amoalu_io_mask = pstore1_mask;
  assign amoalu_io_cmd = pstore1_cmd;
  assign amoalu_io_lhs = {s2_data_corrected_hi,s2_data_corrected_lo};
  assign amoalu_io_rhs = pstore1_data;
  assign tag_array_RW0_en = s0_clk_en | _T_19;
  assign tag_array_RW0_wmode = metaArb_io_out_bits_write;
  assign tag_array_RW0_addr = metaArb_io_out_bits_idx;
  always @(posedge tlb_clock) begin
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_7) begin
            tlb_sectored_entries_0_0_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_7) begin
            tlb_sectored_entries_0_0_data_0 <= tlb__GEN_61;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_7) begin
            tlb_sectored_entries_0_0_data_1 <= tlb__GEN_62;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_7) begin
            tlb_sectored_entries_0_0_data_2 <= tlb__GEN_63;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_7) begin
            tlb_sectored_entries_0_0_data_3 <= tlb__GEN_64;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_0_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_174) begin
          tlb_sectored_entries_0_0_valid_0 <= tlb__GEN_669;
        end else begin
          tlb_sectored_entries_0_0_valid_0 <= tlb__GEN_665;
        end
      end else begin
        tlb_sectored_entries_0_0_valid_0 <= tlb__GEN_685;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_0_valid_0 <= tlb__GEN_289;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_0_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_174) begin
          tlb_sectored_entries_0_0_valid_1 <= tlb__GEN_670;
        end else begin
          tlb_sectored_entries_0_0_valid_1 <= tlb__GEN_666;
        end
      end else begin
        tlb_sectored_entries_0_0_valid_1 <= tlb__GEN_686;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_0_valid_1 <= tlb__GEN_290;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_0_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_174) begin
          tlb_sectored_entries_0_0_valid_2 <= tlb__GEN_671;
        end else begin
          tlb_sectored_entries_0_0_valid_2 <= tlb__GEN_667;
        end
      end else begin
        tlb_sectored_entries_0_0_valid_2 <= tlb__GEN_687;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_0_valid_2 <= tlb__GEN_291;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_0_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_174) begin
          tlb_sectored_entries_0_0_valid_3 <= tlb__GEN_672;
        end else begin
          tlb_sectored_entries_0_0_valid_3 <= tlb__GEN_668;
        end
      end else begin
        tlb_sectored_entries_0_0_valid_3 <= tlb__GEN_688;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_0_valid_3 <= tlb__GEN_292;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_9) begin
            tlb_sectored_entries_0_1_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_9) begin
            tlb_sectored_entries_0_1_data_0 <= tlb__GEN_88;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_9) begin
            tlb_sectored_entries_0_1_data_1 <= tlb__GEN_89;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_9) begin
            tlb_sectored_entries_0_1_data_2 <= tlb__GEN_90;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_9) begin
            tlb_sectored_entries_0_1_data_3 <= tlb__GEN_91;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_1_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_579) begin
          tlb_sectored_entries_0_1_valid_0 <= tlb__GEN_701;
        end else begin
          tlb_sectored_entries_0_1_valid_0 <= tlb__GEN_697;
        end
      end else begin
        tlb_sectored_entries_0_1_valid_0 <= tlb__GEN_717;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_1_valid_0 <= tlb__GEN_300;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_1_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_579) begin
          tlb_sectored_entries_0_1_valid_1 <= tlb__GEN_702;
        end else begin
          tlb_sectored_entries_0_1_valid_1 <= tlb__GEN_698;
        end
      end else begin
        tlb_sectored_entries_0_1_valid_1 <= tlb__GEN_718;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_1_valid_1 <= tlb__GEN_301;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_1_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_579) begin
          tlb_sectored_entries_0_1_valid_2 <= tlb__GEN_703;
        end else begin
          tlb_sectored_entries_0_1_valid_2 <= tlb__GEN_699;
        end
      end else begin
        tlb_sectored_entries_0_1_valid_2 <= tlb__GEN_719;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_1_valid_2 <= tlb__GEN_302;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_1_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_579) begin
          tlb_sectored_entries_0_1_valid_3 <= tlb__GEN_704;
        end else begin
          tlb_sectored_entries_0_1_valid_3 <= tlb__GEN_700;
        end
      end else begin
        tlb_sectored_entries_0_1_valid_3 <= tlb__GEN_720;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_1_valid_3 <= tlb__GEN_303;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_11) begin
            tlb_sectored_entries_0_2_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_11) begin
            tlb_sectored_entries_0_2_data_0 <= tlb__GEN_115;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_11) begin
            tlb_sectored_entries_0_2_data_1 <= tlb__GEN_116;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_11) begin
            tlb_sectored_entries_0_2_data_2 <= tlb__GEN_117;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_11) begin
            tlb_sectored_entries_0_2_data_3 <= tlb__GEN_118;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_2_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_984) begin
          tlb_sectored_entries_0_2_valid_0 <= tlb__GEN_733;
        end else begin
          tlb_sectored_entries_0_2_valid_0 <= tlb__GEN_729;
        end
      end else begin
        tlb_sectored_entries_0_2_valid_0 <= tlb__GEN_749;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_2_valid_0 <= tlb__GEN_311;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_2_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_984) begin
          tlb_sectored_entries_0_2_valid_1 <= tlb__GEN_734;
        end else begin
          tlb_sectored_entries_0_2_valid_1 <= tlb__GEN_730;
        end
      end else begin
        tlb_sectored_entries_0_2_valid_1 <= tlb__GEN_750;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_2_valid_1 <= tlb__GEN_312;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_2_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_984) begin
          tlb_sectored_entries_0_2_valid_2 <= tlb__GEN_735;
        end else begin
          tlb_sectored_entries_0_2_valid_2 <= tlb__GEN_731;
        end
      end else begin
        tlb_sectored_entries_0_2_valid_2 <= tlb__GEN_751;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_2_valid_2 <= tlb__GEN_313;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_2_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_984) begin
          tlb_sectored_entries_0_2_valid_3 <= tlb__GEN_736;
        end else begin
          tlb_sectored_entries_0_2_valid_3 <= tlb__GEN_732;
        end
      end else begin
        tlb_sectored_entries_0_2_valid_3 <= tlb__GEN_752;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_2_valid_3 <= tlb__GEN_314;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_13) begin
            tlb_sectored_entries_0_3_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_13) begin
            tlb_sectored_entries_0_3_data_0 <= tlb__GEN_142;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_13) begin
            tlb_sectored_entries_0_3_data_1 <= tlb__GEN_143;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_13) begin
            tlb_sectored_entries_0_3_data_2 <= tlb__GEN_144;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_13) begin
            tlb_sectored_entries_0_3_data_3 <= tlb__GEN_145;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_3_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1389) begin
          tlb_sectored_entries_0_3_valid_0 <= tlb__GEN_765;
        end else begin
          tlb_sectored_entries_0_3_valid_0 <= tlb__GEN_761;
        end
      end else begin
        tlb_sectored_entries_0_3_valid_0 <= tlb__GEN_781;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_3_valid_0 <= tlb__GEN_322;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_3_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1389) begin
          tlb_sectored_entries_0_3_valid_1 <= tlb__GEN_766;
        end else begin
          tlb_sectored_entries_0_3_valid_1 <= tlb__GEN_762;
        end
      end else begin
        tlb_sectored_entries_0_3_valid_1 <= tlb__GEN_782;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_3_valid_1 <= tlb__GEN_323;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_3_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1389) begin
          tlb_sectored_entries_0_3_valid_2 <= tlb__GEN_767;
        end else begin
          tlb_sectored_entries_0_3_valid_2 <= tlb__GEN_763;
        end
      end else begin
        tlb_sectored_entries_0_3_valid_2 <= tlb__GEN_783;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_3_valid_2 <= tlb__GEN_324;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_3_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1389) begin
          tlb_sectored_entries_0_3_valid_3 <= tlb__GEN_768;
        end else begin
          tlb_sectored_entries_0_3_valid_3 <= tlb__GEN_764;
        end
      end else begin
        tlb_sectored_entries_0_3_valid_3 <= tlb__GEN_784;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_3_valid_3 <= tlb__GEN_325;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_15) begin
            tlb_sectored_entries_0_4_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_15) begin
            tlb_sectored_entries_0_4_data_0 <= tlb__GEN_169;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_15) begin
            tlb_sectored_entries_0_4_data_1 <= tlb__GEN_170;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_15) begin
            tlb_sectored_entries_0_4_data_2 <= tlb__GEN_171;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_15) begin
            tlb_sectored_entries_0_4_data_3 <= tlb__GEN_172;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_4_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1794) begin
          tlb_sectored_entries_0_4_valid_0 <= tlb__GEN_797;
        end else begin
          tlb_sectored_entries_0_4_valid_0 <= tlb__GEN_793;
        end
      end else begin
        tlb_sectored_entries_0_4_valid_0 <= tlb__GEN_813;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_4_valid_0 <= tlb__GEN_333;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_4_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1794) begin
          tlb_sectored_entries_0_4_valid_1 <= tlb__GEN_798;
        end else begin
          tlb_sectored_entries_0_4_valid_1 <= tlb__GEN_794;
        end
      end else begin
        tlb_sectored_entries_0_4_valid_1 <= tlb__GEN_814;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_4_valid_1 <= tlb__GEN_334;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_4_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1794) begin
          tlb_sectored_entries_0_4_valid_2 <= tlb__GEN_799;
        end else begin
          tlb_sectored_entries_0_4_valid_2 <= tlb__GEN_795;
        end
      end else begin
        tlb_sectored_entries_0_4_valid_2 <= tlb__GEN_815;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_4_valid_2 <= tlb__GEN_335;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_4_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_1794) begin
          tlb_sectored_entries_0_4_valid_3 <= tlb__GEN_800;
        end else begin
          tlb_sectored_entries_0_4_valid_3 <= tlb__GEN_796;
        end
      end else begin
        tlb_sectored_entries_0_4_valid_3 <= tlb__GEN_816;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_4_valid_3 <= tlb__GEN_336;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_17) begin
            tlb_sectored_entries_0_5_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_17) begin
            tlb_sectored_entries_0_5_data_0 <= tlb__GEN_196;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_17) begin
            tlb_sectored_entries_0_5_data_1 <= tlb__GEN_197;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_17) begin
            tlb_sectored_entries_0_5_data_2 <= tlb__GEN_198;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_17) begin
            tlb_sectored_entries_0_5_data_3 <= tlb__GEN_199;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_5_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2199) begin
          tlb_sectored_entries_0_5_valid_0 <= tlb__GEN_829;
        end else begin
          tlb_sectored_entries_0_5_valid_0 <= tlb__GEN_825;
        end
      end else begin
        tlb_sectored_entries_0_5_valid_0 <= tlb__GEN_845;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_5_valid_0 <= tlb__GEN_344;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_5_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2199) begin
          tlb_sectored_entries_0_5_valid_1 <= tlb__GEN_830;
        end else begin
          tlb_sectored_entries_0_5_valid_1 <= tlb__GEN_826;
        end
      end else begin
        tlb_sectored_entries_0_5_valid_1 <= tlb__GEN_846;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_5_valid_1 <= tlb__GEN_345;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_5_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2199) begin
          tlb_sectored_entries_0_5_valid_2 <= tlb__GEN_831;
        end else begin
          tlb_sectored_entries_0_5_valid_2 <= tlb__GEN_827;
        end
      end else begin
        tlb_sectored_entries_0_5_valid_2 <= tlb__GEN_847;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_5_valid_2 <= tlb__GEN_346;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_5_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2199) begin
          tlb_sectored_entries_0_5_valid_3 <= tlb__GEN_832;
        end else begin
          tlb_sectored_entries_0_5_valid_3 <= tlb__GEN_828;
        end
      end else begin
        tlb_sectored_entries_0_5_valid_3 <= tlb__GEN_848;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_5_valid_3 <= tlb__GEN_347;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_19) begin
            tlb_sectored_entries_0_6_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_19) begin
            tlb_sectored_entries_0_6_data_0 <= tlb__GEN_223;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_19) begin
            tlb_sectored_entries_0_6_data_1 <= tlb__GEN_224;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_19) begin
            tlb_sectored_entries_0_6_data_2 <= tlb__GEN_225;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_19) begin
            tlb_sectored_entries_0_6_data_3 <= tlb__GEN_226;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_6_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2604) begin
          tlb_sectored_entries_0_6_valid_0 <= tlb__GEN_861;
        end else begin
          tlb_sectored_entries_0_6_valid_0 <= tlb__GEN_857;
        end
      end else begin
        tlb_sectored_entries_0_6_valid_0 <= tlb__GEN_877;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_6_valid_0 <= tlb__GEN_355;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_6_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2604) begin
          tlb_sectored_entries_0_6_valid_1 <= tlb__GEN_862;
        end else begin
          tlb_sectored_entries_0_6_valid_1 <= tlb__GEN_858;
        end
      end else begin
        tlb_sectored_entries_0_6_valid_1 <= tlb__GEN_878;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_6_valid_1 <= tlb__GEN_356;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_6_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2604) begin
          tlb_sectored_entries_0_6_valid_2 <= tlb__GEN_863;
        end else begin
          tlb_sectored_entries_0_6_valid_2 <= tlb__GEN_859;
        end
      end else begin
        tlb_sectored_entries_0_6_valid_2 <= tlb__GEN_879;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_6_valid_2 <= tlb__GEN_357;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_6_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_2604) begin
          tlb_sectored_entries_0_6_valid_3 <= tlb__GEN_864;
        end else begin
          tlb_sectored_entries_0_6_valid_3 <= tlb__GEN_860;
        end
      end else begin
        tlb_sectored_entries_0_6_valid_3 <= tlb__GEN_880;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_6_valid_3 <= tlb__GEN_358;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_21) begin
            tlb_sectored_entries_0_7_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_21) begin
            tlb_sectored_entries_0_7_data_0 <= tlb__GEN_250;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_21) begin
            tlb_sectored_entries_0_7_data_1 <= tlb__GEN_251;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_21) begin
            tlb_sectored_entries_0_7_data_2 <= tlb__GEN_252;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (!(tlb__T_2)) begin
          if (tlb__T_21) begin
            tlb_sectored_entries_0_7_data_3 <= tlb__GEN_253;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_7_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3009) begin
          tlb_sectored_entries_0_7_valid_0 <= tlb__GEN_893;
        end else begin
          tlb_sectored_entries_0_7_valid_0 <= tlb__GEN_889;
        end
      end else begin
        tlb_sectored_entries_0_7_valid_0 <= tlb__GEN_909;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_7_valid_0 <= tlb__GEN_366;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_7_valid_1 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3009) begin
          tlb_sectored_entries_0_7_valid_1 <= tlb__GEN_894;
        end else begin
          tlb_sectored_entries_0_7_valid_1 <= tlb__GEN_890;
        end
      end else begin
        tlb_sectored_entries_0_7_valid_1 <= tlb__GEN_910;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_7_valid_1 <= tlb__GEN_367;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_7_valid_2 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3009) begin
          tlb_sectored_entries_0_7_valid_2 <= tlb__GEN_895;
        end else begin
          tlb_sectored_entries_0_7_valid_2 <= tlb__GEN_891;
        end
      end else begin
        tlb_sectored_entries_0_7_valid_2 <= tlb__GEN_911;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_7_valid_2 <= tlb__GEN_368;
      end
    end
    if (tlb__T_4470) begin
      tlb_sectored_entries_0_7_valid_3 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__T_3009) begin
          tlb_sectored_entries_0_7_valid_3 <= tlb__GEN_896;
        end else begin
          tlb_sectored_entries_0_7_valid_3 <= tlb__GEN_892;
        end
      end else begin
        tlb_sectored_entries_0_7_valid_3 <= tlb__GEN_912;
      end
    end else if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        tlb_sectored_entries_0_7_valid_3 <= tlb__GEN_369;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_3) begin
            tlb_superpage_entries_0_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_3) begin
            tlb_superpage_entries_0_data_0 <= tlb__special_entry_data_0_T;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_superpage_entries_0_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__superpage_hits_T_4) begin
          tlb_superpage_entries_0_valid_0 <= 1'h0;
        end else begin
          tlb_superpage_entries_0_valid_0 <= tlb__GEN_498;
        end
      end else begin
        tlb_superpage_entries_0_valid_0 <= tlb__GEN_920;
      end
    end else begin
      tlb_superpage_entries_0_valid_0 <= tlb__GEN_498;
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_4) begin
            tlb_superpage_entries_1_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_4) begin
            tlb_superpage_entries_1_data_0 <= tlb__special_entry_data_0_T;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_superpage_entries_1_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__superpage_hits_T_13) begin
          tlb_superpage_entries_1_valid_0 <= 1'h0;
        end else begin
          tlb_superpage_entries_1_valid_0 <= tlb__GEN_503;
        end
      end else begin
        tlb_superpage_entries_1_valid_0 <= tlb__GEN_925;
      end
    end else begin
      tlb_superpage_entries_1_valid_0 <= tlb__GEN_503;
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_5) begin
            tlb_superpage_entries_2_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_5) begin
            tlb_superpage_entries_2_data_0 <= tlb__special_entry_data_0_T;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_superpage_entries_2_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__superpage_hits_T_22) begin
          tlb_superpage_entries_2_valid_0 <= 1'h0;
        end else begin
          tlb_superpage_entries_2_valid_0 <= tlb__GEN_508;
        end
      end else begin
        tlb_superpage_entries_2_valid_0 <= tlb__GEN_930;
      end
    end else begin
      tlb_superpage_entries_2_valid_0 <= tlb__GEN_508;
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_6) begin
            tlb_superpage_entries_3_tag_vpn <= tlb_r_refill_tag;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (!(tlb__T)) begin
        if (tlb__T_2) begin
          if (tlb__T_6) begin
            tlb_superpage_entries_3_data_0 <= tlb__special_entry_data_0_T;
          end
        end
      end
    end
    if (tlb__T_4470) begin
      tlb_superpage_entries_3_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__superpage_hits_T_31) begin
          tlb_superpage_entries_3_valid_0 <= 1'h0;
        end else begin
          tlb_superpage_entries_3_valid_0 <= tlb__GEN_513;
        end
      end else begin
        tlb_superpage_entries_3_valid_0 <= tlb__GEN_935;
      end
    end else begin
      tlb_superpage_entries_3_valid_0 <= tlb__GEN_513;
    end
    if (tlb_io_ptw_resp_valid) begin
      if (tlb__T) begin
        tlb_special_entry_level <= tlb_io_ptw_resp_bits_level;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (tlb__T) begin
        tlb_special_entry_tag_vpn <= tlb_r_refill_tag;
      end
    end
    if (tlb_io_ptw_resp_valid) begin
      if (tlb__T) begin
        tlb_special_entry_data_0 <= tlb__special_entry_data_0_T;
      end
    end
    if (tlb__T_4470) begin
      tlb_special_entry_valid_0 <= 1'h0;
    end else if (tlb_io_sfence_valid) begin
      if (tlb_io_sfence_bits_rs1) begin
        if (tlb__hitsVec_T_97) begin
          tlb_special_entry_valid_0 <= 1'h0;
        end else begin
          tlb_special_entry_valid_0 <= tlb__GEN_493;
        end
      end else begin
        tlb_special_entry_valid_0 <= tlb__GEN_940;
      end
    end else begin
      tlb_special_entry_valid_0 <= tlb__GEN_493;
    end
    if (tlb_reset) begin
      tlb_state <= 2'h0;
    end else if (tlb_io_ptw_resp_valid) begin
      tlb_state <= 2'h0;
    end else if (tlb__T_53) begin
      tlb_state <= 2'h3;
    end else if (tlb__invalidate_refill_T) begin
      tlb_state <= tlb__GEN_656;
    end else begin
      tlb_state <= tlb__GEN_644;
    end
    if (tlb__T_50) begin
      tlb_r_refill_tag <= tlb_vpn;
    end
    if (tlb__T_50) begin
      if (tlb__r_superpage_repl_addr_T_4) begin
        tlb_r_superpage_repl_addr <= tlb__r_superpage_repl_addr_T_3;
      end else if (tlb__r_superpage_repl_addr_T_6) begin
        tlb_r_superpage_repl_addr <= 2'h0;
      end else if (tlb__r_superpage_repl_addr_T_7) begin
        tlb_r_superpage_repl_addr <= 2'h1;
      end else begin
        tlb_r_superpage_repl_addr <= tlb__r_superpage_repl_addr_T_10;
      end
    end
    if (tlb__T_50) begin
      if (tlb__r_sectored_repl_addr_T_10) begin
        tlb_r_sectored_repl_addr <= tlb__r_sectored_repl_addr_T_9;
      end else if (tlb__r_sectored_repl_addr_T_12) begin
        tlb_r_sectored_repl_addr <= 3'h0;
      end else if (tlb__r_sectored_repl_addr_T_13) begin
        tlb_r_sectored_repl_addr <= 3'h1;
      end else begin
        tlb_r_sectored_repl_addr <= tlb__r_sectored_repl_addr_T_24;
      end
    end
    if (tlb__T_50) begin
      tlb_r_sectored_hit_valid <= tlb__T_30;
    end
    if (tlb__T_50) begin
      tlb_r_sectored_hit_bits <= tlb__T_38;
    end
    if (tlb__T_50) begin
      tlb_r_need_gpa <= tlb_tlb_hit_if_not_gpa_miss;
    end
    if (tlb_reset) begin
      tlb_state_vec_0 <= 7'h0;
    end else if (tlb__T_23) begin
      if (tlb__T_30) begin
        tlb_state_vec_0 <= tlb__state_vec_0_T_22;
      end
    end
    if (tlb_reset) begin
      tlb_state_reg_1 <= 3'h0;
    end else if (tlb__T_23) begin
      if (tlb__T_41) begin
        tlb_state_reg_1 <= tlb__state_reg_T_8;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (tlb__T_60 & (tlb_io_sfence_valid & tlb__T_59)) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (tlb_io_sfence_valid & tlb__T_59 & tlb__T_60) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TLB.scala:486 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= s1_valid_x12;
    end
    if (reset) begin
      lrscCount <= 7'h0;
    end else if (s1_probe) begin
      lrscCount <= 7'h0;
    end else if (s2_valid_masked & lrscValid) begin
      lrscCount <= 7'h3;
    end else if (_lrscBackingOff_T) begin
      lrscCount <= _lrscCount_T_2;
    end else begin
      lrscCount <= _GEN_143;
    end
    if (reset) begin
      s1_probe <= 1'h0;
    end else begin
      s1_probe <= _GEN_323;
    end
    if (reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    if (reset) begin
      release_state <= 4'h0;
    end else if (_T_337) begin
      release_state <= 4'h0;
    end else if (_T_333) begin
      if (releaseDone) begin
        release_state <= 4'h6;
      end else begin
        release_state <= _GEN_345;
      end
    end else begin
      release_state <= _GEN_345;
    end
    if (reset) begin
      release_ack_wait <= 1'h0;
    end else if (_T_333) begin
      release_ack_wait <= _GEN_354;
    end else if (_T_292) begin
      if (!(grantIsCached)) begin
        release_ack_wait <= _GEN_228;
      end
    end
    if (_T_333) begin
      if (_T_318 & c_first) begin
        release_ack_addr <= probe_bits_address;
      end
    end
    if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s2_valid_x44;
    end
    if (s2_want_victimize) begin
      probe_bits_address <= res_2_address;
    end
    if (s1_probe) begin
      s2_probe_state_state <= s1_meta_hit_state_state;
    end
    if (reset) begin
      counter_1 <= 10'h0;
    end else if (_T_318) begin
      if (c_first) begin
        if (beats1_opdata_1) begin
          counter_1 <= beats1_decode_1;
        end else begin
          counter_1 <= 10'h0;
        end
      end else begin
        counter_1 <= counter1_1;
      end
    end
    s2_release_data_valid <= s1_release_data_valid & ~releaseRejected;
    if (s0_clk_en) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (_T_292) begin
      if (grantIsCached) begin
        s2_req_cmd <= _GEN_65;
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_cmd <= 5'h0;
        end else begin
          s2_req_cmd <= _GEN_65;
        end
      end else begin
        s2_req_cmd <= _GEN_65;
      end
    end else begin
      s2_req_cmd <= _GEN_65;
    end
    if (reset) begin
      pstore1_held <= 1'h0;
    end else begin
      pstore1_held <= pstore1_valid & pstore2_valid & ~pstore_drain;
    end
    if (_pstore1_cmd_T) begin
      pstore1_addr <= s1_vaddr;
    end
    if (s0_clk_en) begin
      s1_req_addr <= s0_req_addr;
    end
    if (_pstore1_cmd_T) begin
      if (_s1_write_T_1) begin
        pstore1_mask <= io_cpu_s1_data_mask;
      end else begin
        pstore1_mask <= s1_mask_xwr;
      end
    end
    if (s0_clk_en) begin
      s1_req_size <= io_cpu_req_bits_size;
    end
    if (reset) begin
      pstore2_valid <= 1'h0;
    end else begin
      pstore2_valid <= pstore2_valid & _pstore1_held_T_9 | advance_pstore1;
    end
    if (advance_pstore1) begin
      pstore2_addr <= pstore1_addr;
    end
    if (advance_pstore1) begin
      mask <= _pstore2_storegen_mask_mask_T_2;
    end
    s2_not_nacked_in_s1 <= ~s1_nack;
    if (_T_74) begin
      s2_hit_state_state <= s1_meta_hit_state_state;
    end
    if (s0_clk_en) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if (s0_clk_en) begin
      s1_req_signed <= io_cpu_req_bits_signed;
    end
    if (s0_clk_en) begin
      s1_req_dprv <= io_cpu_req_bits_dprv;
    end
    if (s0_clk_en) begin
      s1_tlb_req_vaddr <= s0_req_addr;
    end
    if (s0_clk_en) begin
      s1_tlb_req_passthrough <= s0_req_phys;
    end
    if (s0_clk_en) begin
      s1_tlb_req_size <= io_cpu_req_bits_size;
    end
    if (s0_clk_en) begin
      s1_tlb_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (s0_clk_en) begin
      s1_tlb_req_prv <= io_cpu_req_bits_dprv;
    end
    s1_flush_valid <= _s1_flush_valid_T & _T_45 & _s2_cannot_victimize_T & _io_cpu_req_ready_T & _tl_out_a_valid_T_7;
    flushed <= reset | _GEN_406;
    if (reset) begin
      flushing <= 1'h0;
    end else if (flushing) begin
      if (flushed & _io_cpu_req_ready_T & _tl_out_a_valid_T_7) begin
        flushing <= 1'h0;
      end else begin
        flushing <= _GEN_386;
      end
    end else begin
      flushing <= _GEN_386;
    end
    if (_T_345) begin
      if (_metaArb_io_in_5_valid_T & _tl_out_a_valid_T_7 & _s2_valid_cached_miss_T_3) begin
        flushing_req_size <= s2_req_size;
      end
    end
    if (reset) begin
      cached_grant_wait <= 1'h0;
    end else if (_T_292) begin
      if (grantIsCached) begin
        if (d_last) begin
          cached_grant_wait <= 1'h0;
        end else begin
          cached_grant_wait <= _GEN_203;
        end
      end else begin
        cached_grant_wait <= _GEN_203;
      end
    end else begin
      cached_grant_wait <= _GEN_203;
    end
    if (reset) begin
      resetting <= 1'h0;
    end else if (resetting) begin
      if (flushDone) begin
        resetting <= 1'h0;
      end else begin
        resetting <= _GEN_372;
      end
    end else begin
      resetting <= _GEN_372;
    end
    if (reset) begin
      flushCounter <= 8'hc0;
    end else begin
      flushCounter <= _GEN_409[7:0];
    end
    if (_T_284) begin
      if (!(s2_uncached)) begin
        if (s2_hit_valid) begin
          refill_way <= s2_hit_way;
        end else begin
          refill_way <= s2_victim_way;
        end
      end
    end
    if (reset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (_T_292) begin
      if (grantIsCached) begin
        uncachedInFlight_0 <= _GEN_190;
      end else if (grantIsUncached) begin
        uncachedInFlight_0 <= _GEN_211;
      end else begin
        uncachedInFlight_0 <= _GEN_190;
      end
    end else begin
      uncachedInFlight_0 <= _GEN_190;
    end
    if (_T_284) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_addr <= s2_req_addr;
        end
      end
    end
    if (_T_284) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_tag <= s2_req_tag;
        end
      end
    end
    if (_T_284) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_size <= s2_req_size;
        end
      end
    end
    if (_T_284) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_signed <= s2_req_signed;
        end
      end
    end
    if (s0_clk_en) begin
      s1_did_read <= _s1_did_read_T_54;
    end
    if (s1_valid_not_nacked) begin
      s2_hit_way <= s1_meta_hit_way;
    end
    if (_T_74) begin
      if (flushing) begin
        s2_victim_way_r <= flushCounter[7:6];
      end else begin
        s2_victim_way_r <= lfsr[1:0];
      end
    end
    if (s1_probe) begin
      s2_probe_way <= s1_meta_hit_way;
    end
    if (_T_292) begin
      if (grantIsCached) begin
        s2_req_addr <= _GEN_63;
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_addr <= _s2_req_addr_T_1;
        end else begin
          s2_req_addr <= _GEN_63;
        end
      end else begin
        s2_req_addr <= _GEN_63;
      end
    end else begin
      s2_req_addr <= _GEN_63;
    end
    if (_T_292) begin
      if (grantIsCached) begin
        s2_req_tag <= _GEN_64;
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_tag <= uncachedReqs_0_tag;
        end else begin
          s2_req_tag <= _GEN_64;
        end
      end else begin
        s2_req_tag <= _GEN_64;
      end
    end else begin
      s2_req_tag <= _GEN_64;
    end
    if (_T_292) begin
      if (grantIsCached) begin
        s2_req_size <= _GEN_66;
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_size <= uncachedReqs_0_size;
        end else begin
          s2_req_size <= _GEN_66;
        end
      end else begin
        s2_req_size <= _GEN_66;
      end
    end else begin
      s2_req_size <= _GEN_66;
    end
    if (_T_292) begin
      if (grantIsCached) begin
        s2_req_signed <= _GEN_67;
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_signed <= uncachedReqs_0_signed;
        end else begin
          s2_req_signed <= _GEN_67;
        end
      end else begin
        s2_req_signed <= _GEN_67;
      end
    end else begin
      s2_req_signed <= _GEN_67;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_req_dprv <= s1_req_dprv;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_tlb_xcpt_pf_ld <= tlb_io_resp_pf_ld;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_tlb_xcpt_pf_st <= tlb_io_resp_pf_st;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_tlb_xcpt_ae_ld <= tlb_io_resp_ae_ld;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_tlb_xcpt_ae_st <= tlb_io_resp_ae_st;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_tlb_xcpt_ma_ld <= tlb_io_resp_ma_ld;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_tlb_xcpt_ma_st <= tlb_io_resp_ma_st;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin
      s2_pma_cacheable <= tlb_io_resp_cacheable;
    end
    if (_T_292) begin
      if (!(grantIsCached)) begin
        if (grantIsUncached) begin
          if (grantIsUncachedData) begin
            s2_uncached_resp_addr <= uncachedReqs_0_addr;
          end
        end
      end
    end
    if (_T_74) begin
      s2_vaddr_r <= s1_vaddr;
    end
    s2_flush_valid_pre_tag_ecc <= s1_flush_valid;
    if (s1_meta_clk_en) begin
      s2_meta_corrected_r <= tag_array_RW0_rdata_0;
    end
    if (s1_meta_clk_en) begin
      s2_meta_corrected_r_1 <= tag_array_RW0_rdata_1;
    end
    if (s1_meta_clk_en) begin
      s2_meta_corrected_r_2 <= tag_array_RW0_rdata_2;
    end
    if (s1_meta_clk_en) begin
      s2_meta_corrected_r_3 <= tag_array_RW0_rdata_3;
    end
    if (grantIsUncachedData & (blockUncachedGrant | s1_valid)) begin
      if (auto_out_d_valid) begin
        blockUncachedGrant <= _T_312;
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid;
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid;
    end
    if (reset) begin
      counter <= 10'h0;
    end else if (_T_292) begin
      if (d_first) begin
        if (beats1_opdata) begin
          counter <= beats1_decode;
        end else begin
          counter <= 10'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (en) begin
      s2_data <= _s2_data_T_15;
    end
    if (s2_valid_hit_pre_data_ecc_and_waw & _c_cat_T_48 & _io_cpu_req_ready_T_1 | s2_valid_cached_miss) begin
      lrscAddr <= s2_req_addr[31:6];
    end
    if (_pstore1_cmd_T) begin
      pstore1_cmd <= s1_req_cmd;
    end
    if (_pstore1_cmd_T) begin
      pstore1_data <= io_cpu_s1_data_data;
    end
    if (_pstore1_cmd_T) begin
      pstore1_way <= s1_meta_hit_way;
    end
    if (_pstore1_cmd_T) begin
      pstore1_rmw_r <= _pstore1_rmw_T_52;
    end
    pstore_drain_on_miss_REG <= io_cpu_s2_nack;
    if (advance_pstore1) begin
      pstore2_way <= pstore1_way;
    end
    if (advance_pstore1) begin
      pstore2_storegen_data_r <= pstore1_storegen_data[7:0];
    end
    if (advance_pstore1) begin
      pstore2_storegen_data_r_1 <= pstore1_storegen_data[15:8];
    end
    if (advance_pstore1) begin
      pstore2_storegen_data_r_2 <= pstore1_storegen_data[23:16];
    end
    if (advance_pstore1) begin
      pstore2_storegen_data_r_3 <= pstore1_storegen_data[31:24];
    end
    s1_release_data_valid <= dataArb_io_in_2_ready & dataArb_io_in_2_valid;
    io_cpu_s2_xcpt_REG <= tlb_io_req_valid & _s1_valid_not_nacked_T;
    doUncachedResp <= io_cpu_replay_next;
    REG <= reset;
    if (reset) begin
      io_cpu_perf_release_counter <= 10'h0;
    end else if (_T_318) begin
      if (io_cpu_perf_release_first) begin
        if (beats1_opdata_1) begin
          io_cpu_perf_release_counter <= beats1_decode_1;
        end else begin
          io_cpu_perf_release_counter <= 10'h0;
        end
      end else begin
        io_cpu_perf_release_counter <= io_cpu_perf_release_counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_dataArb_io_in_3_valid_T_52 | res) & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_dataArb_io_in_3_valid_T_52 | res)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1158 assert(!needsRead(req) || res)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(s1_valid_masked & _s1_write_T_1) | &_T_68) & _dataArb_io_in_3_valid_T_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_dataArb_io_in_3_valid_T_56 & ~(~(s1_valid_masked & _s1_write_T_1) | &_T_68)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:302 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_dataArb_io_in_3_valid_T_52 | res) & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_dataArb_io_in_3_valid_T_52 | res)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1158 assert(!needsRead(req) || res)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(pstore1_rmw_r | _T_275 == pstore1_valid) & _dataArb_io_in_3_valid_T_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_dataArb_io_in_3_valid_T_56 & ~(pstore1_rmw_r | _T_275 == pstore1_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:483 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_io_cpu_req_ready_T_1 & (_T_292 & grantIsCached & _dataArb_io_in_3_valid_T_56)) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_292 & grantIsCached & _dataArb_io_in_3_valid_T_56 & _io_cpu_req_ready_T_1) begin
          $fwrite(32'h80000002,
            "Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:650 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_a_source_T & (_T_292 & _T_369 & grantIsUncached & _T_297 & _dataArb_io_in_3_valid_T_56)) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_292 & _T_369 & grantIsUncached & _T_297 & _dataArb_io_in_3_valid_T_56 & _a_source_T) begin
          $fwrite(32'h80000002,
            "Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:660 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_tl_out_a_valid_T_7 & (_GEN_481 & _tl_d_data_encoded_T_8 & grantIsVoluntary & _dataArb_io_in_3_valid_T_56)
          ) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_481 & _tl_d_data_encoded_T_8 & grantIsVoluntary & _dataArb_io_in_3_valid_T_56 & _tl_out_a_valid_T_7
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:681 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_304 == (_T_292 & d_first & grantIsCached)) & _dataArb_io_in_3_valid_T_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_dataArb_io_in_3_valid_T_56 & ~(_T_304 == (_T_292 & d_first & grantIsCached))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:689 assert(tl_out.e.fire() === (tl_out.d.fire() && d_first && grantIsCached))\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(s2_valid_flush_line | s2_flush_valid_pre_tag_ecc | io_cpu_s2_nack) & (s2_want_victimize &
          _dataArb_io_in_3_valid_T_56)) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_want_victimize & _dataArb_io_in_3_valid_T_56 & ~(s2_valid_flush_line | s2_flush_valid_pre_tag_ecc |
          io_cpu_s2_nack)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:790 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n"
            );
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_io_cpu_s2_nack_T_4 & (doUncachedResp & _dataArb_io_in_3_valid_T_56)) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & _dataArb_io_in_3_valid_T_56 & ~_io_cpu_s2_nack_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:924 assert(!s2_valid_hit)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_sectored_entries_0_0_tag_vpn = _RAND_0[19:0];
  _RAND_1 = {2{`RANDOM}};
  tlb_sectored_entries_0_0_data_0 = _RAND_1[40:0];
  _RAND_2 = {2{`RANDOM}};
  tlb_sectored_entries_0_0_data_1 = _RAND_2[40:0];
  _RAND_3 = {2{`RANDOM}};
  tlb_sectored_entries_0_0_data_2 = _RAND_3[40:0];
  _RAND_4 = {2{`RANDOM}};
  tlb_sectored_entries_0_0_data_3 = _RAND_4[40:0];
  _RAND_5 = {1{`RANDOM}};
  tlb_sectored_entries_0_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tlb_sectored_entries_0_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  tlb_sectored_entries_0_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tlb_sectored_entries_0_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  tlb_sectored_entries_0_1_tag_vpn = _RAND_9[19:0];
  _RAND_10 = {2{`RANDOM}};
  tlb_sectored_entries_0_1_data_0 = _RAND_10[40:0];
  _RAND_11 = {2{`RANDOM}};
  tlb_sectored_entries_0_1_data_1 = _RAND_11[40:0];
  _RAND_12 = {2{`RANDOM}};
  tlb_sectored_entries_0_1_data_2 = _RAND_12[40:0];
  _RAND_13 = {2{`RANDOM}};
  tlb_sectored_entries_0_1_data_3 = _RAND_13[40:0];
  _RAND_14 = {1{`RANDOM}};
  tlb_sectored_entries_0_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  tlb_sectored_entries_0_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  tlb_sectored_entries_0_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tlb_sectored_entries_0_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  tlb_sectored_entries_0_2_tag_vpn = _RAND_18[19:0];
  _RAND_19 = {2{`RANDOM}};
  tlb_sectored_entries_0_2_data_0 = _RAND_19[40:0];
  _RAND_20 = {2{`RANDOM}};
  tlb_sectored_entries_0_2_data_1 = _RAND_20[40:0];
  _RAND_21 = {2{`RANDOM}};
  tlb_sectored_entries_0_2_data_2 = _RAND_21[40:0];
  _RAND_22 = {2{`RANDOM}};
  tlb_sectored_entries_0_2_data_3 = _RAND_22[40:0];
  _RAND_23 = {1{`RANDOM}};
  tlb_sectored_entries_0_2_valid_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  tlb_sectored_entries_0_2_valid_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  tlb_sectored_entries_0_2_valid_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tlb_sectored_entries_0_2_valid_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  tlb_sectored_entries_0_3_tag_vpn = _RAND_27[19:0];
  _RAND_28 = {2{`RANDOM}};
  tlb_sectored_entries_0_3_data_0 = _RAND_28[40:0];
  _RAND_29 = {2{`RANDOM}};
  tlb_sectored_entries_0_3_data_1 = _RAND_29[40:0];
  _RAND_30 = {2{`RANDOM}};
  tlb_sectored_entries_0_3_data_2 = _RAND_30[40:0];
  _RAND_31 = {2{`RANDOM}};
  tlb_sectored_entries_0_3_data_3 = _RAND_31[40:0];
  _RAND_32 = {1{`RANDOM}};
  tlb_sectored_entries_0_3_valid_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tlb_sectored_entries_0_3_valid_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tlb_sectored_entries_0_3_valid_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tlb_sectored_entries_0_3_valid_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tlb_sectored_entries_0_4_tag_vpn = _RAND_36[19:0];
  _RAND_37 = {2{`RANDOM}};
  tlb_sectored_entries_0_4_data_0 = _RAND_37[40:0];
  _RAND_38 = {2{`RANDOM}};
  tlb_sectored_entries_0_4_data_1 = _RAND_38[40:0];
  _RAND_39 = {2{`RANDOM}};
  tlb_sectored_entries_0_4_data_2 = _RAND_39[40:0];
  _RAND_40 = {2{`RANDOM}};
  tlb_sectored_entries_0_4_data_3 = _RAND_40[40:0];
  _RAND_41 = {1{`RANDOM}};
  tlb_sectored_entries_0_4_valid_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  tlb_sectored_entries_0_4_valid_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  tlb_sectored_entries_0_4_valid_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tlb_sectored_entries_0_4_valid_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  tlb_sectored_entries_0_5_tag_vpn = _RAND_45[19:0];
  _RAND_46 = {2{`RANDOM}};
  tlb_sectored_entries_0_5_data_0 = _RAND_46[40:0];
  _RAND_47 = {2{`RANDOM}};
  tlb_sectored_entries_0_5_data_1 = _RAND_47[40:0];
  _RAND_48 = {2{`RANDOM}};
  tlb_sectored_entries_0_5_data_2 = _RAND_48[40:0];
  _RAND_49 = {2{`RANDOM}};
  tlb_sectored_entries_0_5_data_3 = _RAND_49[40:0];
  _RAND_50 = {1{`RANDOM}};
  tlb_sectored_entries_0_5_valid_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  tlb_sectored_entries_0_5_valid_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  tlb_sectored_entries_0_5_valid_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  tlb_sectored_entries_0_5_valid_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  tlb_sectored_entries_0_6_tag_vpn = _RAND_54[19:0];
  _RAND_55 = {2{`RANDOM}};
  tlb_sectored_entries_0_6_data_0 = _RAND_55[40:0];
  _RAND_56 = {2{`RANDOM}};
  tlb_sectored_entries_0_6_data_1 = _RAND_56[40:0];
  _RAND_57 = {2{`RANDOM}};
  tlb_sectored_entries_0_6_data_2 = _RAND_57[40:0];
  _RAND_58 = {2{`RANDOM}};
  tlb_sectored_entries_0_6_data_3 = _RAND_58[40:0];
  _RAND_59 = {1{`RANDOM}};
  tlb_sectored_entries_0_6_valid_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  tlb_sectored_entries_0_6_valid_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  tlb_sectored_entries_0_6_valid_2 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  tlb_sectored_entries_0_6_valid_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  tlb_sectored_entries_0_7_tag_vpn = _RAND_63[19:0];
  _RAND_64 = {2{`RANDOM}};
  tlb_sectored_entries_0_7_data_0 = _RAND_64[40:0];
  _RAND_65 = {2{`RANDOM}};
  tlb_sectored_entries_0_7_data_1 = _RAND_65[40:0];
  _RAND_66 = {2{`RANDOM}};
  tlb_sectored_entries_0_7_data_2 = _RAND_66[40:0];
  _RAND_67 = {2{`RANDOM}};
  tlb_sectored_entries_0_7_data_3 = _RAND_67[40:0];
  _RAND_68 = {1{`RANDOM}};
  tlb_sectored_entries_0_7_valid_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  tlb_sectored_entries_0_7_valid_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  tlb_sectored_entries_0_7_valid_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  tlb_sectored_entries_0_7_valid_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  tlb_superpage_entries_0_tag_vpn = _RAND_72[19:0];
  _RAND_73 = {2{`RANDOM}};
  tlb_superpage_entries_0_data_0 = _RAND_73[40:0];
  _RAND_74 = {1{`RANDOM}};
  tlb_superpage_entries_0_valid_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  tlb_superpage_entries_1_tag_vpn = _RAND_75[19:0];
  _RAND_76 = {2{`RANDOM}};
  tlb_superpage_entries_1_data_0 = _RAND_76[40:0];
  _RAND_77 = {1{`RANDOM}};
  tlb_superpage_entries_1_valid_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  tlb_superpage_entries_2_tag_vpn = _RAND_78[19:0];
  _RAND_79 = {2{`RANDOM}};
  tlb_superpage_entries_2_data_0 = _RAND_79[40:0];
  _RAND_80 = {1{`RANDOM}};
  tlb_superpage_entries_2_valid_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  tlb_superpage_entries_3_tag_vpn = _RAND_81[19:0];
  _RAND_82 = {2{`RANDOM}};
  tlb_superpage_entries_3_data_0 = _RAND_82[40:0];
  _RAND_83 = {1{`RANDOM}};
  tlb_superpage_entries_3_valid_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  tlb_special_entry_level = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  tlb_special_entry_tag_vpn = _RAND_85[19:0];
  _RAND_86 = {2{`RANDOM}};
  tlb_special_entry_data_0 = _RAND_86[40:0];
  _RAND_87 = {1{`RANDOM}};
  tlb_special_entry_valid_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  tlb_state = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  tlb_r_refill_tag = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  tlb_r_superpage_repl_addr = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  tlb_r_sectored_repl_addr = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  tlb_r_sectored_hit_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  tlb_r_sectored_hit_bits = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  tlb_r_need_gpa = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  tlb_state_vec_0 = _RAND_95[6:0];
  _RAND_96 = {1{`RANDOM}};
  tlb_state_reg_1 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  s1_valid = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lrscCount = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  s1_probe = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  s2_probe = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  release_state = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  release_ack_wait = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  release_ack_addr = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  s2_valid = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  probe_bits_address = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  s2_probe_state_state = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  counter_1 = _RAND_107[9:0];
  _RAND_108 = {1{`RANDOM}};
  s2_release_data_valid = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  s1_req_cmd = _RAND_109[4:0];
  _RAND_110 = {1{`RANDOM}};
  s2_req_cmd = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  pstore1_held = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  pstore1_addr = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  s1_req_addr = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  pstore1_mask = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  s1_req_size = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  pstore2_valid = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  pstore2_addr = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mask = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  s2_not_nacked_in_s1 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  s2_hit_state_state = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  s1_req_tag = _RAND_121[6:0];
  _RAND_122 = {1{`RANDOM}};
  s1_req_signed = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  s1_req_dprv = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  s1_tlb_req_vaddr = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  s1_tlb_req_passthrough = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  s1_tlb_req_size = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  s1_tlb_req_cmd = _RAND_127[4:0];
  _RAND_128 = {1{`RANDOM}};
  s1_tlb_req_prv = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  s1_flush_valid = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  flushed = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  flushing = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  flushing_req_size = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  cached_grant_wait = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  resetting = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  flushCounter = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  refill_way = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  uncachedInFlight_0 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  uncachedReqs_0_addr = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  uncachedReqs_0_tag = _RAND_139[6:0];
  _RAND_140 = {1{`RANDOM}};
  uncachedReqs_0_size = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  uncachedReqs_0_signed = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  s1_did_read = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  s2_hit_way = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  s2_victim_way_r = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  s2_probe_way = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  s2_req_addr = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  s2_req_tag = _RAND_147[6:0];
  _RAND_148 = {1{`RANDOM}};
  s2_req_size = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  s2_req_signed = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  s2_req_dprv = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_ld = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_st = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_ld = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_st = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_ld = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_st = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  s2_pma_cacheable = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  s2_uncached_resp_addr = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  s2_vaddr_r = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  s2_flush_valid_pre_tag_ecc = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  s2_meta_corrected_r = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  s2_meta_corrected_r_1 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  s2_meta_corrected_r_2 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  s2_meta_corrected_r_3 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  blockUncachedGrant = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  counter = _RAND_166[9:0];
  _RAND_167 = {1{`RANDOM}};
  s2_data = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  lrscAddr = _RAND_168[25:0];
  _RAND_169 = {1{`RANDOM}};
  pstore1_cmd = _RAND_169[4:0];
  _RAND_170 = {1{`RANDOM}};
  pstore1_data = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  pstore1_way = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  pstore1_rmw_r = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  pstore_drain_on_miss_REG = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  pstore2_way = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  pstore2_storegen_data_r = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  pstore2_storegen_data_r_1 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  pstore2_storegen_data_r_2 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  pstore2_storegen_data_r_3 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  s1_release_data_valid = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  io_cpu_s2_xcpt_REG = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  doUncachedResp = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  REG = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  io_cpu_perf_release_counter = _RAND_183[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule