// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef __ERVP_PLATFORM_CONTROLLER_MEMORYMAP_OFFSET_H__
`define __ERVP_PLATFORM_CONTROLLER_MEMORYMAP_OFFSET_H__

`define BW_MMAP_OFFSET_ERVP_PLATFORM_CONTROLLER 18
`define ERVP_PLATFORM_CONTROLLER_ADDR_INTERVAL 8
`define BW_UNUSED_ERVP_PLATFORM_CONTROLLER 3
`define NUM_ERVP_PLATFORM_CONTROLLER_SUBMODULE 4
`define BW_SEL_ERVP_PLATFORM_CONTROLLER_SUBMODULE 2
`define SUBMODULE_INDEX_ERVP_PLATFORM_CONTROLLER_RESET 0
`define SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_RESET (32'h 0)
`define SUBMODULE_INDEX_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER 1
`define SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER (32'h 10000)
`define SUBMODULE_INDEX_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO 2
`define SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO (32'h 20000)
`define SUBMODULE_INDEX_ERVP_PLATFORM_CONTROLLER_EXTERNAL 3
`define SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_EXTERNAL (32'h 30000)

`define BW_MMAP_SUBOFFSET_RESET 5
`define BW_UNUSED_RESET 3
`define MMAP_SUBOFFSET_RESET_CMD (32'h 0)
`define MMAP_SUBOFFSET_RESET_MASK (32'h 8)
`define MMAP_SUBOFFSET_RESET_SEQUENCE (32'h 10)

`define MMAP_OFFSET_RESET_CMD (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_RESET+`MMAP_SUBOFFSET_RESET_CMD)
`define MMAP_OFFSET_RESET_MASK (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_RESET+`MMAP_SUBOFFSET_RESET_MASK)
`define MMAP_OFFSET_RESET_SEQUENCE (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_RESET+`MMAP_SUBOFFSET_RESET_SEQUENCE)

`define BW_MMAP_SUBOFFSET_PLATFORM_REGISTER 8
`define BW_UNUSED_PLATFORM_REGISTER 3
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_BOOT_MODE (32'h 0)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_INITIALIZED (32'h 8)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_SIM_ENV (32'h 10)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_JTAG_SELECT (32'h 18)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_BOOT_STATUS (32'h 20)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_APP_ADDR (32'h 28)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_PROC_AUTO_ID (32'h 30)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_PROC_STATUS (32'h 38)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC00 (32'h 40)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC01 (32'h 48)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC02 (32'h 50)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC03 (32'h 58)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST00 (32'h 60)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST01 (32'h 68)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST02 (32'h 70)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST03 (32'h 78)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_IMP_TYPE (32'h 80)
`define MMAP_SUBOFFSET_PLATFORM_REGISTER_FLASH_BASE_ADDR (32'h 88)

`define MMAP_OFFSET_PLATFORM_REGISTER_BOOT_MODE (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_BOOT_MODE)
`define MMAP_OFFSET_PLATFORM_REGISTER_INITIALIZED (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_INITIALIZED)
`define MMAP_OFFSET_PLATFORM_REGISTER_SIM_ENV (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_SIM_ENV)
`define MMAP_OFFSET_PLATFORM_REGISTER_JTAG_SELECT (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_JTAG_SELECT)
`define MMAP_OFFSET_PLATFORM_REGISTER_BOOT_STATUS (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_BOOT_STATUS)
`define MMAP_OFFSET_PLATFORM_REGISTER_APP_ADDR (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_APP_ADDR)
`define MMAP_OFFSET_PLATFORM_REGISTER_PROC_AUTO_ID (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_PROC_AUTO_ID)
`define MMAP_OFFSET_PLATFORM_REGISTER_PROC_STATUS (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_PROC_STATUS)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_PC00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC00)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_PC01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC01)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_PC02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC02)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_PC03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_PC03)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_INST00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST00)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_INST01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST01)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_INST02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST02)
`define MMAP_OFFSET_PLATFORM_REGISTER_CORE_INST03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_CORE_INST03)
`define MMAP_OFFSET_PLATFORM_REGISTER_IMP_TYPE (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_IMP_TYPE)
`define MMAP_OFFSET_PLATFORM_REGISTER_FLASH_BASE_ADDR (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_PLATFORM_REGISTER+`MMAP_SUBOFFSET_PLATFORM_REGISTER_FLASH_BASE_ADDR)

`define BW_MMAP_SUBOFFSET_DESIGN_INFO 8
`define BW_UNUSED_DESIGN_INFO 3
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE00 (32'h 0)
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE01 (32'h 8)
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE02 (32'h 10)
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE03 (32'h 18)
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE04 (32'h 20)
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE05 (32'h 28)
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE06 (32'h 30)
`define MMAP_SUBOFFSET_DESIGN_INFO_DATE07 (32'h 38)
`define MMAP_SUBOFFSET_DESIGN_INFO_USERNAME00 (32'h 40)
`define MMAP_SUBOFFSET_DESIGN_INFO_USERNAME01 (32'h 48)
`define MMAP_SUBOFFSET_DESIGN_INFO_USERNAME02 (32'h 50)
`define MMAP_SUBOFFSET_DESIGN_INFO_USERNAME03 (32'h 58)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME00 (32'h 60)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME01 (32'h 68)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME02 (32'h 70)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME03 (32'h 78)
`define MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME00 (32'h 80)
`define MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME01 (32'h 88)
`define MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME02 (32'h 90)
`define MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME03 (32'h 98)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION00 (32'h a0)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION01 (32'h a8)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION02 (32'h b0)
`define MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION03 (32'h b8)
`define MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION00 (32'h c0)
`define MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION01 (32'h c8)
`define MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION02 (32'h d0)
`define MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION03 (32'h d8)

`define MMAP_OFFSET_DESIGN_INFO_DATE00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE00)
`define MMAP_OFFSET_DESIGN_INFO_DATE01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE01)
`define MMAP_OFFSET_DESIGN_INFO_DATE02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE02)
`define MMAP_OFFSET_DESIGN_INFO_DATE03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE03)
`define MMAP_OFFSET_DESIGN_INFO_DATE04 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE04)
`define MMAP_OFFSET_DESIGN_INFO_DATE05 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE05)
`define MMAP_OFFSET_DESIGN_INFO_DATE06 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE06)
`define MMAP_OFFSET_DESIGN_INFO_DATE07 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DATE07)
`define MMAP_OFFSET_DESIGN_INFO_USERNAME00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_USERNAME00)
`define MMAP_OFFSET_DESIGN_INFO_USERNAME01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_USERNAME01)
`define MMAP_OFFSET_DESIGN_INFO_USERNAME02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_USERNAME02)
`define MMAP_OFFSET_DESIGN_INFO_USERNAME03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_USERNAME03)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_NAME00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME00)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_NAME01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME01)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_NAME02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME02)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_NAME03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_NAME03)
`define MMAP_OFFSET_DESIGN_INFO_PLATFORM_NAME00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME00)
`define MMAP_OFFSET_DESIGN_INFO_PLATFORM_NAME01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME01)
`define MMAP_OFFSET_DESIGN_INFO_PLATFORM_NAME02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME02)
`define MMAP_OFFSET_DESIGN_INFO_PLATFORM_NAME03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_PLATFORM_NAME03)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_VERSION00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION00)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_VERSION01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION01)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_VERSION02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION02)
`define MMAP_OFFSET_DESIGN_INFO_HOME_GIT_VERSION03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_HOME_GIT_VERSION03)
`define MMAP_OFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION00 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION00)
`define MMAP_OFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION01 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION01)
`define MMAP_OFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION02 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION02)
`define MMAP_OFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION03 (`SUBMODULE_ADDR_ERVP_PLATFORM_CONTROLLER_DESIGN_INFO+`MMAP_SUBOFFSET_DESIGN_INFO_DEVKIT_GIT_VERSION03)

`define BW_MMAP_SUBOFFSET_EXTERNAL 16
`define BW_UNUSED_EXTERNAL 3

`define BW_RESET_CMD 3
`define RESET_CMD_DEFAULT_VALUE 0
`define RESET_CMD_IDLE 0
`define RESET_CMD_INIT 1
`define RESET_CMD_AUTO_INCR 2
`define RESET_CMD_NEXT_STEP 3
`define RESET_CMD_IDLE_WITH_ERROR 4
`define RESET_CMD_INDEX_INIT 0
`define RESET_CMD_INDEX_AUTO_INCR 1
`define RESET_CMD_INDEX_IDLE_WITH_ERROR 2

`define BW_RESET_MASK 32
`define RESET_MASK_DEFAULT_VALUE 0

`define BW_RESET_SEQUENCE 32
`define RESET_SEQUENCE_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_BOOT_MODE 4
`define PLATFORM_REGISTER_BOOT_MODE_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_INITIALIZED 1
`define PLATFORM_REGISTER_INITIALIZED_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_SIM_ENV 1
`define PLATFORM_REGISTER_SIM_ENV_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_JTAG_SELECT 1
`define PLATFORM_REGISTER_JTAG_SELECT_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_BOOT_STATUS 32
`define PLATFORM_REGISTER_BOOT_STATUS_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_APP_ADDR 32
`define PLATFORM_REGISTER_APP_ADDR_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_PROC_AUTO_ID 32
`define PLATFORM_REGISTER_PROC_AUTO_ID_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_PROC_STATUS 32
`define PLATFORM_REGISTER_PROC_STATUS_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_CORE_PC 32
`define PLATFORM_REGISTER_CORE_PC_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_CORE_INST 32
`define PLATFORM_REGISTER_CORE_INST_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_IMP_TYPE 32
`define PLATFORM_REGISTER_IMP_TYPE_DEFAULT_VALUE 0

`define BW_PLATFORM_REGISTER_FLASH_BASE_ADDR 32
`define PLATFORM_REGISTER_FLASH_BASE_ADDR_DEFAULT_VALUE 0

`define BW_DESIGN_INFO_DATE 32
`define DESIGN_INFO_DATE_DEFAULT_VALUE 0

`define BW_DESIGN_INFO_USERNAME 32
`define DESIGN_INFO_USERNAME_DEFAULT_VALUE 0

`define BW_DESIGN_INFO_HOME_GIT_NAME 32
`define DESIGN_INFO_HOME_GIT_NAME_DEFAULT_VALUE 0

`define BW_DESIGN_INFO_PLATFORM_NAME 32
`define DESIGN_INFO_PLATFORM_NAME_DEFAULT_VALUE 0

`define BW_DESIGN_INFO_HOME_GIT_VERSION 32
`define DESIGN_INFO_HOME_GIT_VERSION_DEFAULT_VALUE 0

`define BW_DESIGN_INFO_DEVKIT_GIT_VERSION 32
`define DESIGN_INFO_DEVKIT_GIT_VERSION_DEFAULT_VALUE 0

`define BW_BOOT_MODE 1
`define BOOT_MODE_DEFAULT_VALUE 0
`define BOOT_MODE_OCD 0
`define BOOT_MODE_STAND_ALONE 1
`define BOOT_MODE_INDEX_STAND_ALONE 0

`define BW_BOOT_STATUS 2
`define BOOT_STATUS_DEFAULT_VALUE 0
`define BOOT_STATUS_RESETED 0
`define BOOT_STATUS_APP_LOAD 1
`define BOOT_STATUS_ALL_READY 2
`define BOOT_STATUS_INDEX_APP_LOAD 0
`define BOOT_STATUS_INDEX_ALL_READY 1

`define BW_JTAG_SELECT 1
`define JTAG_SELECT_DEFAULT_VALUE 0
`define JTAG_SELECT_NOC 0
`define JTAG_SELECT_CORE 1
`define JTAG_SELECT_INDEX_CORE 0

`define BW_IMP_TYPE 2
`define IMP_TYPE_DEFAULT_VALUE 0
`define IMP_TYPE_RTL 0
`define IMP_TYPE_FPGA 1
`define IMP_TYPE_CHIP 2
`define IMP_TYPE_VP 3
`define IMP_TYPE_INDEX_FPGA 0
`define IMP_TYPE_INDEX_CHIP 1

`endif