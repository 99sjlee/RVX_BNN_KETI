// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_019
`define RVX_GDEF_019

`define RVX_GDEF_297 5
`define RVX_GDEF_076 8
`define RVX_GDEF_251 3
`define RVX_GDEF_092 1

`define RVX_GDEF_008 (32'h 0)
`define RVX_GDEF_095 (32'h 8)
`define RVX_GDEF_181 (32'h 10)

`define RVX_GDEF_091 (`RVX_GDEF_008)
`define RVX_GDEF_054 (`RVX_GDEF_095)
`define RVX_GDEF_105 (`RVX_GDEF_181)

`define RVX_GDEF_355 32
`define RVX_GDEF_193 0

`define RVX_GDEF_239 32
`define RVX_GDEF_332 0

`define RVX_GDEF_209 2
`define RVX_GDEF_314 0

`define RVX_GDEF_139 5
`define RVX_GDEF_393 0
`define RVX_GDEF_166 1
`define RVX_GDEF_331 2
`define RVX_GDEF_308 4
`define RVX_GDEF_226 8
`define RVX_GDEF_403 16
`define RVX_GDEF_361 0
`define RVX_GDEF_271 1
`define RVX_GDEF_132 2
`define RVX_GDEF_027 3
`define RVX_GDEF_320 4
`define RVX_GDEF_376 0

`define RVX_GDEF_408 2
`define RVX_GDEF_245 0
`define RVX_GDEF_196 0
`define RVX_GDEF_404 1
`define RVX_GDEF_385 2
`define RVX_GDEF_034 3
`define RVX_GDEF_045 0
`define RVX_GDEF_270 1

`define RVX_GDEF_089 3
`define RVX_GDEF_136 0
`define RVX_GDEF_156 0
`define RVX_GDEF_023 1
`define RVX_GDEF_369 2
`define RVX_GDEF_189 3
`define RVX_GDEF_290 4
`define RVX_GDEF_295 5
`define RVX_GDEF_211 0
`define RVX_GDEF_016 1
`define RVX_GDEF_366 2

`endif