// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_231
`define RVX_GDEF_231

`define RVX_GDEF_028 None
`define RVX_GDEF_021 8
`define RVX_GDEF_282 3
`define RVX_GDEF_219 0

`define RVX_GDEF_053 5
`define RVX_GDEF_073 0
`define RVX_GDEF_155 0
`define RVX_GDEF_125 16
`define RVX_GDEF_407 20
`define RVX_GDEF_301 21
`define RVX_GDEF_059 22
`define RVX_GDEF_421 23
`define RVX_GDEF_035 24
`define RVX_GDEF_382 28

`define RVX_GDEF_372 5
`define RVX_GDEF_427 0
`define RVX_GDEF_379 16
`define RVX_GDEF_396 4
`define RVX_GDEF_164 1
`define RVX_GDEF_224 1
`define RVX_GDEF_094 1
`define RVX_GDEF_395 1
`define RVX_GDEF_176 1
`define RVX_GDEF_162 3

`endif