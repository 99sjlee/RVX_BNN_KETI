// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_261
`define RVX_GDEF_261

`define RVX_GDEF_082 8
`define RVX_GDEF_323 8
`define RVX_GDEF_174 3
`define RVX_GDEF_266 1

`define RVX_GDEF_328 (32'h 0)
`define RVX_GDEF_391 (32'h 8)
`define RVX_GDEF_099 (32'h 10)
`define RVX_GDEF_128 (32'h 18)
`define RVX_GDEF_030 (32'h 20)
`define RVX_GDEF_252 (32'h 28)
`define RVX_GDEF_191 (32'h 30)
`define RVX_GDEF_052 (32'h 38)
`define RVX_GDEF_217 (32'h 40)
`define RVX_GDEF_386 (32'h 48)
`define RVX_GDEF_263 (32'h 50)
`define RVX_GDEF_036 (32'h 58)
`define RVX_GDEF_357 (32'h 60)
`define RVX_GDEF_397 (32'h 68)
`define RVX_GDEF_227 (32'h 70)
`define RVX_GDEF_228 (32'h 78)
`define RVX_GDEF_056 (32'h 80)
`define RVX_GDEF_063 (32'h 88)
`define RVX_GDEF_242 (32'h 90)
`define RVX_GDEF_426 (32'h 98)
`define RVX_GDEF_339 (32'h a0)
`define RVX_GDEF_318 (32'h a8)
`define RVX_GDEF_006 (32'h b0)
`define RVX_GDEF_292 (32'h b8)
`define RVX_GDEF_351 (32'h c0)

`define RVX_GDEF_240 (`RVX_GDEF_328)
`define RVX_GDEF_300 (`RVX_GDEF_391)
`define RVX_GDEF_409 (`RVX_GDEF_099)
`define RVX_GDEF_293 (`RVX_GDEF_128)
`define RVX_GDEF_145 (`RVX_GDEF_030)
`define RVX_GDEF_269 (`RVX_GDEF_252)
`define RVX_GDEF_345 (`RVX_GDEF_191)
`define RVX_GDEF_354 (`RVX_GDEF_052)
`define RVX_GDEF_121 (`RVX_GDEF_217)
`define RVX_GDEF_163 (`RVX_GDEF_386)
`define RVX_GDEF_000 (`RVX_GDEF_263)
`define RVX_GDEF_024 (`RVX_GDEF_036)
`define RVX_GDEF_316 (`RVX_GDEF_357)
`define RVX_GDEF_364 (`RVX_GDEF_397)
`define RVX_GDEF_122 (`RVX_GDEF_227)
`define RVX_GDEF_140 (`RVX_GDEF_228)
`define RVX_GDEF_398 (`RVX_GDEF_056)
`define RVX_GDEF_142 (`RVX_GDEF_063)
`define RVX_GDEF_353 (`RVX_GDEF_242)
`define RVX_GDEF_255 (`RVX_GDEF_426)
`define RVX_GDEF_327 (`RVX_GDEF_339)
`define RVX_GDEF_259 (`RVX_GDEF_318)
`define RVX_GDEF_406 (`RVX_GDEF_006)
`define RVX_GDEF_237 (`RVX_GDEF_292)
`define RVX_GDEF_072 (`RVX_GDEF_351)

`define RVX_GDEF_311 8
`define RVX_GDEF_287 0

`define RVX_GDEF_347 32
`define RVX_GDEF_321 0

`define RVX_GDEF_405 32
`define RVX_GDEF_313 0

`define RVX_GDEF_138 32
`define RVX_GDEF_304 0

`endif