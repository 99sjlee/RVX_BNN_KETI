// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_129
`define RVX_GDEF_129

`define RVX_GDEF_186 15
`define RVX_GDEF_068 8
`define RVX_GDEF_203 3
`define RVX_GDEF_026 5
`define RVX_GDEF_011 3
`define RVX_GDEF_388 0
`define RVX_GDEF_220 (32'h 0)
`define RVX_GDEF_350 1
`define RVX_GDEF_065 (32'h 1000)
`define RVX_GDEF_336 2
`define RVX_GDEF_279 (32'h 2000)
`define RVX_GDEF_365 3
`define RVX_GDEF_088 (32'h 3000)
`define RVX_GDEF_235 4
`define RVX_GDEF_344 (32'h 4000)

`define RVX_GDEF_415 12
`define RVX_GDEF_080 3

`define RVX_GDEF_194 12
`define RVX_GDEF_070 3

`define RVX_GDEF_411 12
`define RVX_GDEF_392 3

`define RVX_GDEF_031 5
`define RVX_GDEF_283 3
`define RVX_GDEF_185 (32'h 0)
`define RVX_GDEF_278 (32'h 8)
`define RVX_GDEF_104 (32'h 10)

`define RVX_GDEF_064 (`RVX_GDEF_088+`RVX_GDEF_185)
`define RVX_GDEF_256 (`RVX_GDEF_088+`RVX_GDEF_278)
`define RVX_GDEF_113 (`RVX_GDEF_088+`RVX_GDEF_104)

`define RVX_GDEF_402 4
`define RVX_GDEF_084 3

`define RVX_GDEF_241 8
`define RVX_GDEF_262 0

`define RVX_GDEF_286 11

`define RVX_GDEF_370 11

`endif