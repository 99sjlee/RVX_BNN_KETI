// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef __ERVP_EXTERNAL_PERI_GROUP_MEMORYMAP_OFFSET_H__
`define __ERVP_EXTERNAL_PERI_GROUP_MEMORYMAP_OFFSET_H__

`define BW_MMAP_OFFSET_ERVP_EXTERNAL_PERI_GROUP 12
`define ERVP_EXTERNAL_PERI_GROUP_ADDR_INTERVAL 8
`define BW_UNUSED_ERVP_EXTERNAL_PERI_GROUP 3
`define NUM_ERVP_EXTERNAL_PERI_GROUP_SUBMODULE 12
`define BW_SEL_ERVP_EXTERNAL_PERI_GROUP_SUBMODULE 4
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC 0
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC (32'h 0)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_UART0 1
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_UART0 (32'h 100)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_UART1 2
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_UART1 (32'h 200)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_UART2 3
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_UART2 (32'h 300)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_UART3 4
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_UART3 (32'h 400)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_I2C0 5
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_I2C0 (32'h 500)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_I2C1 6
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_I2C1 (32'h 600)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_I2C2 7
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_I2C2 (32'h 700)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_I2C3 8
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_I2C3 (32'h 800)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_SPI 9
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPI (32'h 900)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_GPIO 10
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO (32'h a00)
`define SUBMODULE_INDEX_ERVP_EXTERNAL_PERI_GROUP_SPIO 11
`define SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO (32'h b00)

`define BW_MMAP_SUBOFFSET_EPG_MISC 7
`define BW_UNUSED_EPG_MISC 3
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG00 (32'h 0)
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG01 (32'h 8)
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG02 (32'h 10)
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG03 (32'h 18)
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG04 (32'h 20)
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG05 (32'h 28)
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG06 (32'h 30)
`define MMAP_SUBOFFSET_EPG_MISC_EXTREG07 (32'h 38)
`define MMAP_SUBOFFSET_EPG_MISC_GPIO_TICK_CFG (32'h 40)

`define MMAP_OFFSET_EPG_MISC_EXTREG00 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG00)
`define MMAP_OFFSET_EPG_MISC_EXTREG01 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG01)
`define MMAP_OFFSET_EPG_MISC_EXTREG02 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG02)
`define MMAP_OFFSET_EPG_MISC_EXTREG03 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG03)
`define MMAP_OFFSET_EPG_MISC_EXTREG04 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG04)
`define MMAP_OFFSET_EPG_MISC_EXTREG05 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG05)
`define MMAP_OFFSET_EPG_MISC_EXTREG06 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG06)
`define MMAP_OFFSET_EPG_MISC_EXTREG07 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_EXTREG07)
`define MMAP_OFFSET_EPG_MISC_GPIO_TICK_CFG (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_EPG_MISC+`MMAP_SUBOFFSET_EPG_MISC_GPIO_TICK_CFG)

`define BW_MMAP_SUBOFFSET_UART0 8
`define BW_UNUSED_UART0 3

`define BW_MMAP_SUBOFFSET_UART1 8
`define BW_UNUSED_UART1 3

`define BW_MMAP_SUBOFFSET_UART2 8
`define BW_UNUSED_UART2 3

`define BW_MMAP_SUBOFFSET_UART3 8
`define BW_UNUSED_UART3 3

`define BW_MMAP_SUBOFFSET_I2C0 8
`define BW_UNUSED_I2C0 3

`define BW_MMAP_SUBOFFSET_I2C1 8
`define BW_UNUSED_I2C1 3

`define BW_MMAP_SUBOFFSET_I2C2 8
`define BW_UNUSED_I2C2 3

`define BW_MMAP_SUBOFFSET_I2C3 8
`define BW_UNUSED_I2C3 3

`define BW_MMAP_SUBOFFSET_SPI 8
`define BW_UNUSED_SPI 3

`define BW_MMAP_SUBOFFSET_GPIO 7
`define BW_UNUSED_GPIO 3
`define MMAP_SUBOFFSET_GPIO_USER_GPIO00 (32'h 0)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO01 (32'h 8)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO02 (32'h 10)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO03 (32'h 18)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO04 (32'h 20)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO05 (32'h 28)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO06 (32'h 30)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO07 (32'h 38)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO08 (32'h 40)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO09 (32'h 48)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO10 (32'h 50)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO11 (32'h 58)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO12 (32'h 60)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO13 (32'h 68)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO14 (32'h 70)
`define MMAP_SUBOFFSET_GPIO_USER_GPIO15 (32'h 78)

`define MMAP_OFFSET_GPIO_USER_GPIO00 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO00)
`define MMAP_OFFSET_GPIO_USER_GPIO01 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO01)
`define MMAP_OFFSET_GPIO_USER_GPIO02 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO02)
`define MMAP_OFFSET_GPIO_USER_GPIO03 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO03)
`define MMAP_OFFSET_GPIO_USER_GPIO04 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO04)
`define MMAP_OFFSET_GPIO_USER_GPIO05 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO05)
`define MMAP_OFFSET_GPIO_USER_GPIO06 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO06)
`define MMAP_OFFSET_GPIO_USER_GPIO07 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO07)
`define MMAP_OFFSET_GPIO_USER_GPIO08 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO08)
`define MMAP_OFFSET_GPIO_USER_GPIO09 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO09)
`define MMAP_OFFSET_GPIO_USER_GPIO10 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO10)
`define MMAP_OFFSET_GPIO_USER_GPIO11 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO11)
`define MMAP_OFFSET_GPIO_USER_GPIO12 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO12)
`define MMAP_OFFSET_GPIO_USER_GPIO13 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO13)
`define MMAP_OFFSET_GPIO_USER_GPIO14 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO14)
`define MMAP_OFFSET_GPIO_USER_GPIO15 (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_GPIO+`MMAP_SUBOFFSET_GPIO_USER_GPIO15)

`define BW_MMAP_SUBOFFSET_SPIO 7
`define BW_UNUSED_SPIO 3
`define MMAP_SUBOFFSET_SPIO_OLED_DCSEL (32'h 0)
`define MMAP_SUBOFFSET_SPIO_OLED_RSTNN (32'h 8)
`define MMAP_SUBOFFSET_SPIO_OLED_VBAT (32'h 10)
`define MMAP_SUBOFFSET_SPIO_OLED_VDD (32'h 18)
`define MMAP_SUBOFFSET_SPIO_WIFI_RSTNN (32'h 20)
`define MMAP_SUBOFFSET_SPIO_WIFI_WP (32'h 28)
`define MMAP_SUBOFFSET_SPIO_WIFI_HIBERNATE (32'h 30)
`define MMAP_SUBOFFSET_SPIO_WIFI_ITR_CLEAR (32'h 38)
`define MMAP_SUBOFFSET_SPIO_WIFI_ITR_PENDING (32'h 40)
`define MMAP_SUBOFFSET_SPIO_SPI_CS_ACTIVE_LOW (32'h 48)
`define MMAP_SUBOFFSET_SPIO_SPI_SELECT (32'h 50)
`define MMAP_SUBOFFSET_SPIO_AIOIF_CONFIG (32'h 58)
`define MMAP_SUBOFFSET_SPIO_SERIAL_COMM_CONTROL (32'h 60)

`define MMAP_OFFSET_SPIO_OLED_DCSEL (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_OLED_DCSEL)
`define MMAP_OFFSET_SPIO_OLED_RSTNN (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_OLED_RSTNN)
`define MMAP_OFFSET_SPIO_OLED_VBAT (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_OLED_VBAT)
`define MMAP_OFFSET_SPIO_OLED_VDD (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_OLED_VDD)
`define MMAP_OFFSET_SPIO_WIFI_RSTNN (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_WIFI_RSTNN)
`define MMAP_OFFSET_SPIO_WIFI_WP (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_WIFI_WP)
`define MMAP_OFFSET_SPIO_WIFI_HIBERNATE (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_WIFI_HIBERNATE)
`define MMAP_OFFSET_SPIO_WIFI_ITR_CLEAR (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_WIFI_ITR_CLEAR)
`define MMAP_OFFSET_SPIO_WIFI_ITR_PENDING (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_WIFI_ITR_PENDING)
`define MMAP_OFFSET_SPIO_SPI_CS_ACTIVE_LOW (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_SPI_CS_ACTIVE_LOW)
`define MMAP_OFFSET_SPIO_SPI_SELECT (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_SPI_SELECT)
`define MMAP_OFFSET_SPIO_AIOIF_CONFIG (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_AIOIF_CONFIG)
`define MMAP_OFFSET_SPIO_SERIAL_COMM_CONTROL (`SUBMODULE_ADDR_ERVP_EXTERNAL_PERI_GROUP_SPIO+`MMAP_SUBOFFSET_SPIO_SERIAL_COMM_CONTROL)

`define BW_SPIO_SPI_CS_ACTIVE_LOW 32
`define SPIO_SPI_CS_ACTIVE_LOW_DEFAULT_VALUE -1

`define BW_SPIO_SERIAL_COMM_CONTROL 4
`define SPIO_SERIAL_COMM_CONTROL_DEFAULT_VALUE 0
`define SPIO_SERIAL_COMM_CONTROL_SPI_CLK_USER_OE 1
`define SPIO_SERIAL_COMM_CONTROL_SPI_CLK_USER_VALUE 2
`define SPIO_SERIAL_COMM_CONTROL_SPI_DQ0_USER_OE 4
`define SPIO_SERIAL_COMM_CONTROL_SPI_DQ0_USER_VALUE 8
`define SPIO_SERIAL_COMM_CONTROL_INDEX_SPI_CLK_USER_OE 0
`define SPIO_SERIAL_COMM_CONTROL_INDEX_SPI_CLK_USER_VALUE 1
`define SPIO_SERIAL_COMM_CONTROL_INDEX_SPI_DQ0_USER_OE 2
`define SPIO_SERIAL_COMM_CONTROL_INDEX_SPI_DQ0_USER_VALUE 3
`define SPIO_SERIAL_COMM_CONTROL_NONE 0

`define BW_EPG_MISC_EXTREG 32
`define EPG_MISC_EXTREG_DEFAULT_VALUE 0

`define BW_EPG_MISC_GPIO_TICK_CFG 16
`define EPG_MISC_GPIO_TICK_CFG_DEFAULT_VALUE 0

`define BW_GPIO_USER_GPIO 32
`define GPIO_USER_GPIO_DEFAULT_VALUE 0

`define BW_SPIO_OLED_DCSEL 1
`define SPIO_OLED_DCSEL_DEFAULT_VALUE 0

`define BW_SPIO_OLED_RSTNN 1
`define SPIO_OLED_RSTNN_DEFAULT_VALUE 0

`define BW_SPIO_OLED_VBAT 1
`define SPIO_OLED_VBAT_DEFAULT_VALUE 0

`define BW_SPIO_OLED_VDD 1
`define SPIO_OLED_VDD_DEFAULT_VALUE 0

`define BW_SPIO_WIFI_RSTNN 1
`define SPIO_WIFI_RSTNN_DEFAULT_VALUE 0

`define BW_SPIO_WIFI_WP 1
`define SPIO_WIFI_WP_DEFAULT_VALUE 0

`define BW_SPIO_WIFI_HIBERNATE 1
`define SPIO_WIFI_HIBERNATE_DEFAULT_VALUE 0

`define BW_SPIO_WIFI_ITR_CLEAR 1
`define SPIO_WIFI_ITR_CLEAR_DEFAULT_VALUE 0

`define BW_SPIO_WIFI_ITR_PENDING 1
`define SPIO_WIFI_ITR_PENDING_DEFAULT_VALUE 0

`define BW_SPIO_SPI_SELECT 32
`define SPIO_SPI_SELECT_DEFAULT_VALUE 0

`define BW_SPIO_AIOIF_CONFIG 32
`define SPIO_AIOIF_CONFIG_DEFAULT_VALUE 0

`define BW_OLED_DC_SEL 1
`define OLED_DC_SEL_DEFAULT_VALUE 0
`define OLED_DC_SEL_COMMAND 0
`define OLED_DC_SEL_DATA 1
`define OLED_DC_SEL_INDEX_DATA 0

`define BW_OCD_FLASH_CMD 3
`define OCD_FLASH_CMD_DEFAULT_VALUE 0
`define OCD_FLASH_CMD_IDLE 0
`define OCD_FLASH_CMD_CHECK 1
`define OCD_FLASH_CMD_ERASE 2
`define OCD_FLASH_CMD_READ 3
`define OCD_FLASH_CMD_WRITE 4
`define OCD_FLASH_CMD_INDEX_CHECK 0
`define OCD_FLASH_CMD_INDEX_ERASE 1
`define OCD_FLASH_CMD_INDEX_WRITE 2

`define BW_BOOT_STATUS 2
`define BOOT_STATUS_DEFAULT_VALUE 0
`define BOOT_STATUS_RESETED 0
`define BOOT_STATUS_APP_LOAD 1
`define BOOT_STATUS_ALL_READY 2
`define BOOT_STATUS_INDEX_APP_LOAD 0
`define BOOT_STATUS_INDEX_ALL_READY 1

`define BW_GPIO_CONFIG 5
`define GPIO_CONFIG_DEFAULT_VALUE 0
`define GPIO_CONFIG_IS_SIGNED_VALUE 1
`define GPIO_CONFIG_IS_OUTPUT_PORT 2
`define GPIO_CONFIG_ITR_ENABLE 4
`define GPIO_CONFIG_DEBOUNCE_ENABLE 8
`define GPIO_CONFIG_USER_IO_SELECT 16
`define GPIO_CONFIG_INDEX_IS_SIGNED_VALUE 0
`define GPIO_CONFIG_INDEX_IS_OUTPUT_PORT 1
`define GPIO_CONFIG_INDEX_ITR_ENABLE 2
`define GPIO_CONFIG_INDEX_DEBOUNCE_ENABLE 3
`define GPIO_CONFIG_INDEX_USER_IO_SELECT 4
`define GPIO_CONFIG_NONE 0

`define BW_GPIO_CMD 4
`define GPIO_CMD_DEFAULT_VALUE 0
`define GPIO_CMD_WE_VALUE 1
`define GPIO_CMD_WE_CONFIG 2
`define GPIO_CMD_WE_ITR_COND 4
`define GPIO_CMD_CLEAR_ITR 8
`define GPIO_CMD_INDEX_WE_VALUE 0
`define GPIO_CMD_INDEX_WE_CONFIG 1
`define GPIO_CMD_INDEX_WE_ITR_COND 2
`define GPIO_CMD_INDEX_CLEAR_ITR 3
`define GPIO_CMD_NONE 0

`define BW_AIOIF_TYPE 4
`define AIOIF_TYPE_DEFAULT_VALUE 0
`define AIOIF_TYPE_GPIO 1
`define AIOIF_TYPE_I2C 2
`define AIOIF_TYPE_SPI 4
`define AIOIF_TYPE_UART 8
`define AIOIF_TYPE_INDEX_GPIO 0
`define AIOIF_TYPE_INDEX_I2C 1
`define AIOIF_TYPE_INDEX_SPI 2
`define AIOIF_TYPE_INDEX_UART 3
`define AIOIF_TYPE_NONE 0

`define BW_GPIO_VALUE 16
`define GPIO_VALUE_DEFAULT_VALUE 0

`endif