wire [BW_USERNAME-1:0] username_string = `FORMAT_STRING("keti1_arx01");
wire [BW_GIT_NAME-1:0] home_git_name_string = `FORMAT_STRING("_keti_bnn_riscv");
wire [BW_GIT_VERSION-1:0] home_git_version_string = `FORMAT_STRING("1fd523f");
wire [BW_GIT_VERSION-1:0] devkit_git_version_string = `FORMAT_STRING("588e415");
wire [BW_DATE-1:0] design_date_string = `FORMAT_STRING("2025-08-05 11:06");