// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-07-15
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef RVX_GDEF_341
`define RVX_GDEF_341

`define RVX_GDEF_015 6
`define RVX_GDEF_394 8
`define RVX_GDEF_048 3
`define RVX_GDEF_250 1

`define RVX_GDEF_020 (32'h 0)
`define RVX_GDEF_389 (32'h 8)
`define RVX_GDEF_081 (32'h 10)
`define RVX_GDEF_432 (32'h 18)
`define RVX_GDEF_157 (32'h 20)
`define RVX_GDEF_116 (32'h 28)
`define RVX_GDEF_144 (32'h 30)
`define RVX_GDEF_014 (32'h 38)

`define RVX_GDEF_390 (`RVX_GDEF_020)
`define RVX_GDEF_173 (`RVX_GDEF_389)
`define RVX_GDEF_221 (`RVX_GDEF_081)
`define RVX_GDEF_348 (`RVX_GDEF_432)
`define RVX_GDEF_362 (`RVX_GDEF_157)
`define RVX_GDEF_180 (`RVX_GDEF_116)
`define RVX_GDEF_007 (`RVX_GDEF_144)
`define RVX_GDEF_085 (`RVX_GDEF_014)

`define RVX_GDEF_195 3
`define RVX_GDEF_423 0
`define RVX_GDEF_223 0
`define RVX_GDEF_097 1
`define RVX_GDEF_087 2
`define RVX_GDEF_197 3
`define RVX_GDEF_178 4
`define RVX_GDEF_383 0
`define RVX_GDEF_218 1
`define RVX_GDEF_384 2

`define RVX_GDEF_111 1
`define RVX_GDEF_110 0

`define RVX_GDEF_243 32
`define RVX_GDEF_428 0

`define RVX_GDEF_009 32
`define RVX_GDEF_273 0

`define RVX_GDEF_127 32
`define RVX_GDEF_010 0

`define RVX_GDEF_338 32
`define RVX_GDEF_340 0

`define RVX_GDEF_326 32
`define RVX_GDEF_077 0

`define RVX_GDEF_274 32
`define RVX_GDEF_260 0

`define RVX_GDEF_120 2
`define RVX_GDEF_103 0
`define RVX_GDEF_090 0
`define RVX_GDEF_119 1
`define RVX_GDEF_018 2
`define RVX_GDEF_244 3
`define RVX_GDEF_214 0
`define RVX_GDEF_387 1

`define RVX_GDEF_367 16
`define RVX_GDEF_098 0

`define RVX_GDEF_425 16
`define RVX_GDEF_044 0

`define RVX_GDEF_143 16
`define RVX_GDEF_152 0

`endif