`default_nettype wire
module RVCExpander(
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc
);
  wire [6:0] io_out_s_opc = |io_in[12:5] ? 7'h13 : 7'h1f;
  wire [4:0] _io_out_s_T_6 = {2'h1,io_in[4:2]};
  wire [29:0] _io_out_s_T_7 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],io_out_s_opc};
  wire [4:0] io_out_s_0_rs3 = io_in[31:27];
  wire [7:0] _io_out_s_T_15 = {io_in[6:5],io_in[12:10],3'h0};
  wire [4:0] _io_out_s_T_17 = {2'h1,io_in[9:7]};
  wire [27:0] _io_out_s_T_20 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7};
  wire [6:0] _io_out_s_T_31 = {io_in[5],io_in[12:10],io_in[6],2'h0};
  wire [26:0] _io_out_s_T_36 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3};
  wire [26:0] _io_out_s_T_52 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h7};
  wire [26:0] _io_out_s_T_74 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h3f};
  wire [27:0] _io_out_s_T_94 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h27};
  wire [26:0] _io_out_s_T_116 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h23};
  wire [26:0] _io_out_s_T_138 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h27};
  wire [6:0] _io_out_s_T_148 = io_in[12] ? 7'h7f : 7'h0;
  wire [11:0] _io_out_s_T_150 = {_io_out_s_T_148,io_in[6:2]};
  wire [31:0] io_out_s_8_bits = {_io_out_s_T_148,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13};
  wire [9:0] _io_out_s_T_161 = io_in[12] ? 10'h3ff : 10'h0;
  wire [20:0] _io_out_s_T_169 = {_io_out_s_T_161,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0
    };
  wire [31:0] io_out_s_9_bits = {_io_out_s_T_169[20],_io_out_s_T_169[10:1],_io_out_s_T_169[11],_io_out_s_T_169[19:12],5'h1
    ,7'h6f};
  wire [31:0] io_out_s_10_bits = {_io_out_s_T_148,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13};
  wire  _io_out_s_opc_T_7 = |_io_out_s_T_150;
  wire [6:0] io_out_s_opc_1 = |_io_out_s_T_150 ? 7'h37 : 7'h3f;
  wire [14:0] _io_out_s_me_T_2 = io_in[12] ? 15'h7fff : 15'h0;
  wire [31:0] _io_out_s_me_T_4 = {_io_out_s_me_T_2,io_in[6:2],12'h0};
  wire [31:0] io_out_s_me_bits = {_io_out_s_me_T_4[31:12],io_in[11:7],io_out_s_opc_1};
  wire [6:0] io_out_s_opc_2 = _io_out_s_opc_T_7 ? 7'h13 : 7'h1f;
  wire [2:0] _io_out_s_T_230 = io_in[12] ? 3'h7 : 3'h0;
  wire [31:0] io_out_s_res_bits = {_io_out_s_T_230,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:
    7],io_out_s_opc_2};
  wire [31:0] io_out_s_11_bits = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_out_s_res_bits : io_out_s_me_bits;
  wire [4:0] io_out_s_11_rd = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_in[11:7] : io_in[11:7];
  wire [4:0] io_out_s_11_rs2 = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? _io_out_s_T_6 : _io_out_s_T_6;
  wire [4:0] io_out_s_11_rs3 = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_out_s_0_rs3 : io_out_s_0_rs3;
  wire [25:0] _io_out_s_T_251 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13};
  wire [30:0] _GEN_0 = {{5'd0}, _io_out_s_T_251};
  wire [30:0] _io_out_s_T_260 = _GEN_0 | 31'h40000000;
  wire [31:0] _io_out_s_T_270 = {_io_out_s_T_148,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13};
  wire [2:0] _io_out_s_funct_T_2 = {io_in[12],io_in[6:5]};
  wire [2:0] _io_out_s_funct_T_4 = _io_out_s_funct_T_2 == 3'h1 ? 3'h4 : 3'h0;
  wire [2:0] _io_out_s_funct_T_6 = _io_out_s_funct_T_2 == 3'h2 ? 3'h6 : _io_out_s_funct_T_4;
  wire [2:0] _io_out_s_funct_T_8 = _io_out_s_funct_T_2 == 3'h3 ? 3'h7 : _io_out_s_funct_T_6;
  wire [2:0] _io_out_s_funct_T_10 = _io_out_s_funct_T_2 == 3'h4 ? 3'h0 : _io_out_s_funct_T_8;
  wire [2:0] _io_out_s_funct_T_12 = _io_out_s_funct_T_2 == 3'h5 ? 3'h0 : _io_out_s_funct_T_10;
  wire [2:0] _io_out_s_funct_T_14 = _io_out_s_funct_T_2 == 3'h6 ? 3'h2 : _io_out_s_funct_T_12;
  wire [2:0] io_out_s_funct = _io_out_s_funct_T_2 == 3'h7 ? 3'h3 : _io_out_s_funct_T_14;
  wire [30:0] io_out_s_sub = io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h0;
  wire [6:0] io_out_s_opc_3 = io_in[12] ? 7'h3b : 7'h33;
  wire [24:0] _io_out_s_T_277 = {2'h1,io_in[4:2],2'h1,io_in[9:7],io_out_s_funct,2'h1,io_in[9:7],io_out_s_opc_3};
  wire [30:0] _GEN_1 = {{6'd0}, _io_out_s_T_277};
  wire [30:0] _io_out_s_T_278 = _GEN_1 | io_out_s_sub;
  wire [30:0] _io_out_s_T_281 = io_in[11:10] == 2'h1 ? _io_out_s_T_260 : {{5'd0}, _io_out_s_T_251};
  wire [31:0] _io_out_s_T_283 = io_in[11:10] == 2'h2 ? _io_out_s_T_270 : {{1'd0}, _io_out_s_T_281};
  wire [31:0] io_out_s_12_bits = io_in[11:10] == 2'h3 ? {{1'd0}, _io_out_s_T_278} : _io_out_s_T_283;
  wire [31:0] io_out_s_13_bits = {_io_out_s_T_169[20],_io_out_s_T_169[10:1],_io_out_s_T_169[11],_io_out_s_T_169[19:12],5'h0
    ,7'h6f};
  wire [4:0] _io_out_s_T_349 = io_in[12] ? 5'h1f : 5'h0;
  wire [12:0] _io_out_s_T_354 = {_io_out_s_T_349,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0};
  wire [31:0] io_out_s_14_bits = {_io_out_s_T_354[12],_io_out_s_T_354[10:5],5'h0,2'h1,io_in[9:7],3'h0,_io_out_s_T_354[4:
    1],_io_out_s_T_354[11],7'h63};
  wire [31:0] io_out_s_15_bits = {_io_out_s_T_354[12],_io_out_s_T_354[10:5],5'h0,2'h1,io_in[9:7],3'h1,_io_out_s_T_354[4:
    1],_io_out_s_T_354[11],7'h63};
  wire  _io_out_s_load_opc_T_1 = |io_in[11:7];
  wire [6:0] io_out_s_load_opc = |io_in[11:7] ? 7'h3 : 7'h1f;
  wire [25:0] _io_out_s_T_438 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13};
  wire [28:0] _io_out_s_T_448 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7};
  wire [27:0] _io_out_s_T_457 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],io_out_s_load_opc};
  wire [27:0] _io_out_s_T_466 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],7'h7};
  wire [24:0] _io_out_s_mv_T_2 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33};
  wire [24:0] _io_out_s_add_T_3 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33};
  wire [24:0] io_out_s_jr = {io_in[6:2],io_in[11:7],3'h0,12'h67};
  wire [24:0] io_out_s_reserved = {io_out_s_jr[24:7],7'h1f};
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_load_opc_T_1 ? io_out_s_jr : io_out_s_reserved;
  wire  _io_out_s_jr_mv_T_1 = |io_in[6:2];
  wire [31:0] io_out_s_mv_bits = {{7'd0}, _io_out_s_mv_T_2};
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2};
  wire [31:0] io_out_s_jr_mv_bits = |io_in[6:2] ? io_out_s_mv_bits : io_out_s_jr_reserved_bits;
  wire [4:0] io_out_s_jr_mv_rd = |io_in[6:2] ? io_in[11:7] : 5'h0;
  wire [4:0] io_out_s_jr_mv_rs1 = |io_in[6:2] ? 5'h0 : io_in[11:7];
  wire [4:0] io_out_s_jr_mv_rs2 = |io_in[6:2] ? io_in[6:2] : io_in[6:2];
  wire [4:0] io_out_s_jr_mv_rs3 = |io_in[6:2] ? io_out_s_0_rs3 : io_out_s_0_rs3;
  wire [24:0] io_out_s_jalr = {io_in[6:2],io_in[11:7],3'h0,12'he7};
  wire [24:0] _io_out_s_ebreak_T_1 = {io_out_s_jr[24:7],7'h73};
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T_1 | 25'h100000;
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_load_opc_T_1 ? io_out_s_jalr : io_out_s_ebreak;
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T_3};
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2};
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits;
  wire [4:0] io_out_s_jalr_add_rd = _io_out_s_jr_mv_T_1 ? io_in[11:7] : 5'h1;
  wire [4:0] io_out_s_jalr_add_rs1 = _io_out_s_jr_mv_T_1 ? io_in[11:7] : io_in[11:7];
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits;
  wire [4:0] io_out_s_20_rd = io_in[12] ? io_out_s_jalr_add_rd : io_out_s_jr_mv_rd;
  wire [4:0] io_out_s_20_rs1 = io_in[12] ? io_out_s_jalr_add_rs1 : io_out_s_jr_mv_rs1;
  wire [4:0] io_out_s_20_rs2 = io_in[12] ? io_out_s_jr_mv_rs2 : io_out_s_jr_mv_rs2;
  wire [4:0] io_out_s_20_rs3 = io_in[12] ? io_out_s_jr_mv_rs3 : io_out_s_jr_mv_rs3;
  wire [8:0] _io_out_s_T_473 = {io_in[9:7],io_in[12:10],3'h0};
  wire [28:0] _io_out_s_T_480 = {_io_out_s_T_473[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_473[4:0],7'h27};
  wire [7:0] _io_out_s_T_486 = {io_in[8:7],io_in[12:9],2'h0};
  wire [27:0] _io_out_s_T_493 = {_io_out_s_T_486[7:5],io_in[6:2],5'h2,3'h2,_io_out_s_T_486[4:0],7'h23};
  wire [27:0] _io_out_s_T_506 = {_io_out_s_T_486[7:5],io_in[6:2],5'h2,3'h2,_io_out_s_T_486[4:0],7'h27};
  wire [4:0] io_out_s_24_rs1 = io_in[19:15];
  wire [4:0] io_out_s_24_rs2 = io_in[24:20];
  wire [4:0] _io_out_T_2 = {io_in[1:0],io_in[15:13]};
  wire [31:0] io_out_s_1_bits = {{4'd0}, _io_out_s_T_20};
  wire [31:0] io_out_s_0_bits = {{2'd0}, _io_out_s_T_7};
  wire [31:0] _io_out_T_4_bits = _io_out_T_2 == 5'h1 ? io_out_s_1_bits : io_out_s_0_bits;
  wire [4:0] _io_out_T_4_rd = _io_out_T_2 == 5'h1 ? _io_out_s_T_6 : _io_out_s_T_6;
  wire [4:0] _io_out_T_4_rs1 = _io_out_T_2 == 5'h1 ? _io_out_s_T_17 : 5'h2;
  wire [4:0] _io_out_T_4_rs3 = _io_out_T_2 == 5'h1 ? io_out_s_0_rs3 : io_out_s_0_rs3;
  wire [31:0] io_out_s_2_bits = {{5'd0}, _io_out_s_T_36};
  wire [31:0] _io_out_T_6_bits = _io_out_T_2 == 5'h2 ? io_out_s_2_bits : _io_out_T_4_bits;
  wire [4:0] _io_out_T_6_rd = _io_out_T_2 == 5'h2 ? _io_out_s_T_6 : _io_out_T_4_rd;
  wire [4:0] _io_out_T_6_rs1 = _io_out_T_2 == 5'h2 ? _io_out_s_T_17 : _io_out_T_4_rs1;
  wire [4:0] _io_out_T_6_rs3 = _io_out_T_2 == 5'h2 ? io_out_s_0_rs3 : _io_out_T_4_rs3;
  wire [31:0] io_out_s_3_bits = {{5'd0}, _io_out_s_T_52};
  wire [31:0] _io_out_T_8_bits = _io_out_T_2 == 5'h3 ? io_out_s_3_bits : _io_out_T_6_bits;
  wire [4:0] _io_out_T_8_rd = _io_out_T_2 == 5'h3 ? _io_out_s_T_6 : _io_out_T_6_rd;
  wire [4:0] _io_out_T_8_rs1 = _io_out_T_2 == 5'h3 ? _io_out_s_T_17 : _io_out_T_6_rs1;
  wire [4:0] _io_out_T_8_rs3 = _io_out_T_2 == 5'h3 ? io_out_s_0_rs3 : _io_out_T_6_rs3;
  wire [31:0] io_out_s_4_bits = {{5'd0}, _io_out_s_T_74};
  wire [31:0] _io_out_T_10_bits = _io_out_T_2 == 5'h4 ? io_out_s_4_bits : _io_out_T_8_bits;
  wire [4:0] _io_out_T_10_rd = _io_out_T_2 == 5'h4 ? _io_out_s_T_6 : _io_out_T_8_rd;
  wire [4:0] _io_out_T_10_rs1 = _io_out_T_2 == 5'h4 ? _io_out_s_T_17 : _io_out_T_8_rs1;
  wire [4:0] _io_out_T_10_rs3 = _io_out_T_2 == 5'h4 ? io_out_s_0_rs3 : _io_out_T_8_rs3;
  wire [31:0] io_out_s_5_bits = {{4'd0}, _io_out_s_T_94};
  wire [31:0] _io_out_T_12_bits = _io_out_T_2 == 5'h5 ? io_out_s_5_bits : _io_out_T_10_bits;
  wire [4:0] _io_out_T_12_rd = _io_out_T_2 == 5'h5 ? _io_out_s_T_6 : _io_out_T_10_rd;
  wire [4:0] _io_out_T_12_rs1 = _io_out_T_2 == 5'h5 ? _io_out_s_T_17 : _io_out_T_10_rs1;
  wire [4:0] _io_out_T_12_rs3 = _io_out_T_2 == 5'h5 ? io_out_s_0_rs3 : _io_out_T_10_rs3;
  wire [31:0] io_out_s_6_bits = {{5'd0}, _io_out_s_T_116};
  wire [31:0] _io_out_T_14_bits = _io_out_T_2 == 5'h6 ? io_out_s_6_bits : _io_out_T_12_bits;
  wire [4:0] _io_out_T_14_rd = _io_out_T_2 == 5'h6 ? _io_out_s_T_6 : _io_out_T_12_rd;
  wire [4:0] _io_out_T_14_rs1 = _io_out_T_2 == 5'h6 ? _io_out_s_T_17 : _io_out_T_12_rs1;
  wire [4:0] _io_out_T_14_rs3 = _io_out_T_2 == 5'h6 ? io_out_s_0_rs3 : _io_out_T_12_rs3;
  wire [31:0] io_out_s_7_bits = {{5'd0}, _io_out_s_T_138};
  wire [31:0] _io_out_T_16_bits = _io_out_T_2 == 5'h7 ? io_out_s_7_bits : _io_out_T_14_bits;
  wire [4:0] _io_out_T_16_rd = _io_out_T_2 == 5'h7 ? _io_out_s_T_6 : _io_out_T_14_rd;
  wire [4:0] _io_out_T_16_rs1 = _io_out_T_2 == 5'h7 ? _io_out_s_T_17 : _io_out_T_14_rs1;
  wire [4:0] _io_out_T_16_rs3 = _io_out_T_2 == 5'h7 ? io_out_s_0_rs3 : _io_out_T_14_rs3;
  wire [31:0] _io_out_T_18_bits = _io_out_T_2 == 5'h8 ? io_out_s_8_bits : _io_out_T_16_bits;
  wire [4:0] _io_out_T_18_rd = _io_out_T_2 == 5'h8 ? io_in[11:7] : _io_out_T_16_rd;
  wire [4:0] _io_out_T_18_rs1 = _io_out_T_2 == 5'h8 ? io_in[11:7] : _io_out_T_16_rs1;
  wire [4:0] _io_out_T_18_rs2 = _io_out_T_2 == 5'h8 ? _io_out_s_T_6 : _io_out_T_16_rd;
  wire [4:0] _io_out_T_18_rs3 = _io_out_T_2 == 5'h8 ? io_out_s_0_rs3 : _io_out_T_16_rs3;
  wire [31:0] _io_out_T_20_bits = _io_out_T_2 == 5'h9 ? io_out_s_9_bits : _io_out_T_18_bits;
  wire [4:0] _io_out_T_20_rd = _io_out_T_2 == 5'h9 ? 5'h1 : _io_out_T_18_rd;
  wire [4:0] _io_out_T_20_rs1 = _io_out_T_2 == 5'h9 ? io_in[11:7] : _io_out_T_18_rs1;
  wire [4:0] _io_out_T_20_rs2 = _io_out_T_2 == 5'h9 ? _io_out_s_T_6 : _io_out_T_18_rs2;
  wire [4:0] _io_out_T_20_rs3 = _io_out_T_2 == 5'h9 ? io_out_s_0_rs3 : _io_out_T_18_rs3;
  wire [31:0] _io_out_T_22_bits = _io_out_T_2 == 5'ha ? io_out_s_10_bits : _io_out_T_20_bits;
  wire [4:0] _io_out_T_22_rd = _io_out_T_2 == 5'ha ? io_in[11:7] : _io_out_T_20_rd;
  wire [4:0] _io_out_T_22_rs1 = _io_out_T_2 == 5'ha ? 5'h0 : _io_out_T_20_rs1;
  wire [4:0] _io_out_T_22_rs2 = _io_out_T_2 == 5'ha ? _io_out_s_T_6 : _io_out_T_20_rs2;
  wire [4:0] _io_out_T_22_rs3 = _io_out_T_2 == 5'ha ? io_out_s_0_rs3 : _io_out_T_20_rs3;
  wire [31:0] _io_out_T_24_bits = _io_out_T_2 == 5'hb ? io_out_s_11_bits : _io_out_T_22_bits;
  wire [4:0] _io_out_T_24_rd = _io_out_T_2 == 5'hb ? io_out_s_11_rd : _io_out_T_22_rd;
  wire [4:0] _io_out_T_24_rs1 = _io_out_T_2 == 5'hb ? io_out_s_11_rd : _io_out_T_22_rs1;
  wire [4:0] _io_out_T_24_rs2 = _io_out_T_2 == 5'hb ? io_out_s_11_rs2 : _io_out_T_22_rs2;
  wire [4:0] _io_out_T_24_rs3 = _io_out_T_2 == 5'hb ? io_out_s_11_rs3 : _io_out_T_22_rs3;
  wire [31:0] _io_out_T_26_bits = _io_out_T_2 == 5'hc ? io_out_s_12_bits : _io_out_T_24_bits;
  wire [4:0] _io_out_T_26_rd = _io_out_T_2 == 5'hc ? _io_out_s_T_17 : _io_out_T_24_rd;
  wire [4:0] _io_out_T_26_rs1 = _io_out_T_2 == 5'hc ? _io_out_s_T_17 : _io_out_T_24_rs1;
  wire [4:0] _io_out_T_26_rs2 = _io_out_T_2 == 5'hc ? _io_out_s_T_6 : _io_out_T_24_rs2;
  wire [4:0] _io_out_T_26_rs3 = _io_out_T_2 == 5'hc ? io_out_s_0_rs3 : _io_out_T_24_rs3;
  wire [31:0] _io_out_T_28_bits = _io_out_T_2 == 5'hd ? io_out_s_13_bits : _io_out_T_26_bits;
  wire [4:0] _io_out_T_28_rd = _io_out_T_2 == 5'hd ? 5'h0 : _io_out_T_26_rd;
  wire [4:0] _io_out_T_28_rs1 = _io_out_T_2 == 5'hd ? _io_out_s_T_17 : _io_out_T_26_rs1;
  wire [4:0] _io_out_T_28_rs2 = _io_out_T_2 == 5'hd ? _io_out_s_T_6 : _io_out_T_26_rs2;
  wire [4:0] _io_out_T_28_rs3 = _io_out_T_2 == 5'hd ? io_out_s_0_rs3 : _io_out_T_26_rs3;
  wire [31:0] _io_out_T_30_bits = _io_out_T_2 == 5'he ? io_out_s_14_bits : _io_out_T_28_bits;
  wire [4:0] _io_out_T_30_rd = _io_out_T_2 == 5'he ? _io_out_s_T_17 : _io_out_T_28_rd;
  wire [4:0] _io_out_T_30_rs1 = _io_out_T_2 == 5'he ? _io_out_s_T_17 : _io_out_T_28_rs1;
  wire [4:0] _io_out_T_30_rs2 = _io_out_T_2 == 5'he ? 5'h0 : _io_out_T_28_rs2;
  wire [4:0] _io_out_T_30_rs3 = _io_out_T_2 == 5'he ? io_out_s_0_rs3 : _io_out_T_28_rs3;
  wire [31:0] _io_out_T_32_bits = _io_out_T_2 == 5'hf ? io_out_s_15_bits : _io_out_T_30_bits;
  wire [4:0] _io_out_T_32_rd = _io_out_T_2 == 5'hf ? 5'h0 : _io_out_T_30_rd;
  wire [4:0] _io_out_T_32_rs1 = _io_out_T_2 == 5'hf ? _io_out_s_T_17 : _io_out_T_30_rs1;
  wire [4:0] _io_out_T_32_rs2 = _io_out_T_2 == 5'hf ? 5'h0 : _io_out_T_30_rs2;
  wire [4:0] _io_out_T_32_rs3 = _io_out_T_2 == 5'hf ? io_out_s_0_rs3 : _io_out_T_30_rs3;
  wire [31:0] io_out_s_16_bits = {{6'd0}, _io_out_s_T_438};
  wire [31:0] _io_out_T_34_bits = _io_out_T_2 == 5'h10 ? io_out_s_16_bits : _io_out_T_32_bits;
  wire [4:0] _io_out_T_34_rd = _io_out_T_2 == 5'h10 ? io_in[11:7] : _io_out_T_32_rd;
  wire [4:0] _io_out_T_34_rs1 = _io_out_T_2 == 5'h10 ? io_in[11:7] : _io_out_T_32_rs1;
  wire [4:0] _io_out_T_34_rs2 = _io_out_T_2 == 5'h10 ? io_in[6:2] : _io_out_T_32_rs2;
  wire [4:0] _io_out_T_34_rs3 = _io_out_T_2 == 5'h10 ? io_out_s_0_rs3 : _io_out_T_32_rs3;
  wire [31:0] io_out_s_17_bits = {{3'd0}, _io_out_s_T_448};
  wire [31:0] _io_out_T_36_bits = _io_out_T_2 == 5'h11 ? io_out_s_17_bits : _io_out_T_34_bits;
  wire [4:0] _io_out_T_36_rd = _io_out_T_2 == 5'h11 ? io_in[11:7] : _io_out_T_34_rd;
  wire [4:0] _io_out_T_36_rs1 = _io_out_T_2 == 5'h11 ? 5'h2 : _io_out_T_34_rs1;
  wire [4:0] _io_out_T_36_rs2 = _io_out_T_2 == 5'h11 ? io_in[6:2] : _io_out_T_34_rs2;
  wire [4:0] _io_out_T_36_rs3 = _io_out_T_2 == 5'h11 ? io_out_s_0_rs3 : _io_out_T_34_rs3;
  wire [31:0] io_out_s_18_bits = {{4'd0}, _io_out_s_T_457};
  wire [31:0] _io_out_T_38_bits = _io_out_T_2 == 5'h12 ? io_out_s_18_bits : _io_out_T_36_bits;
  wire [4:0] _io_out_T_38_rd = _io_out_T_2 == 5'h12 ? io_in[11:7] : _io_out_T_36_rd;
  wire [4:0] _io_out_T_38_rs1 = _io_out_T_2 == 5'h12 ? 5'h2 : _io_out_T_36_rs1;
  wire [4:0] _io_out_T_38_rs2 = _io_out_T_2 == 5'h12 ? io_in[6:2] : _io_out_T_36_rs2;
  wire [4:0] _io_out_T_38_rs3 = _io_out_T_2 == 5'h12 ? io_out_s_0_rs3 : _io_out_T_36_rs3;
  wire [31:0] io_out_s_19_bits = {{4'd0}, _io_out_s_T_466};
  wire [31:0] _io_out_T_40_bits = _io_out_T_2 == 5'h13 ? io_out_s_19_bits : _io_out_T_38_bits;
  wire [4:0] _io_out_T_40_rd = _io_out_T_2 == 5'h13 ? io_in[11:7] : _io_out_T_38_rd;
  wire [4:0] _io_out_T_40_rs1 = _io_out_T_2 == 5'h13 ? 5'h2 : _io_out_T_38_rs1;
  wire [4:0] _io_out_T_40_rs2 = _io_out_T_2 == 5'h13 ? io_in[6:2] : _io_out_T_38_rs2;
  wire [4:0] _io_out_T_40_rs3 = _io_out_T_2 == 5'h13 ? io_out_s_0_rs3 : _io_out_T_38_rs3;
  wire [31:0] _io_out_T_42_bits = _io_out_T_2 == 5'h14 ? io_out_s_20_bits : _io_out_T_40_bits;
  wire [4:0] _io_out_T_42_rd = _io_out_T_2 == 5'h14 ? io_out_s_20_rd : _io_out_T_40_rd;
  wire [4:0] _io_out_T_42_rs1 = _io_out_T_2 == 5'h14 ? io_out_s_20_rs1 : _io_out_T_40_rs1;
  wire [4:0] _io_out_T_42_rs2 = _io_out_T_2 == 5'h14 ? io_out_s_20_rs2 : _io_out_T_40_rs2;
  wire [4:0] _io_out_T_42_rs3 = _io_out_T_2 == 5'h14 ? io_out_s_20_rs3 : _io_out_T_40_rs3;
  wire [31:0] io_out_s_21_bits = {{3'd0}, _io_out_s_T_480};
  wire [31:0] _io_out_T_44_bits = _io_out_T_2 == 5'h15 ? io_out_s_21_bits : _io_out_T_42_bits;
  wire [4:0] _io_out_T_44_rd = _io_out_T_2 == 5'h15 ? io_in[11:7] : _io_out_T_42_rd;
  wire [4:0] _io_out_T_44_rs1 = _io_out_T_2 == 5'h15 ? 5'h2 : _io_out_T_42_rs1;
  wire [4:0] _io_out_T_44_rs2 = _io_out_T_2 == 5'h15 ? io_in[6:2] : _io_out_T_42_rs2;
  wire [4:0] _io_out_T_44_rs3 = _io_out_T_2 == 5'h15 ? io_out_s_0_rs3 : _io_out_T_42_rs3;
  wire [31:0] io_out_s_22_bits = {{4'd0}, _io_out_s_T_493};
  wire [31:0] _io_out_T_46_bits = _io_out_T_2 == 5'h16 ? io_out_s_22_bits : _io_out_T_44_bits;
  wire [4:0] _io_out_T_46_rd = _io_out_T_2 == 5'h16 ? io_in[11:7] : _io_out_T_44_rd;
  wire [4:0] _io_out_T_46_rs1 = _io_out_T_2 == 5'h16 ? 5'h2 : _io_out_T_44_rs1;
  wire [4:0] _io_out_T_46_rs2 = _io_out_T_2 == 5'h16 ? io_in[6:2] : _io_out_T_44_rs2;
  wire [4:0] _io_out_T_46_rs3 = _io_out_T_2 == 5'h16 ? io_out_s_0_rs3 : _io_out_T_44_rs3;
  wire [31:0] io_out_s_23_bits = {{4'd0}, _io_out_s_T_506};
  wire [31:0] _io_out_T_48_bits = _io_out_T_2 == 5'h17 ? io_out_s_23_bits : _io_out_T_46_bits;
  wire [4:0] _io_out_T_48_rd = _io_out_T_2 == 5'h17 ? io_in[11:7] : _io_out_T_46_rd;
  wire [4:0] _io_out_T_48_rs1 = _io_out_T_2 == 5'h17 ? 5'h2 : _io_out_T_46_rs1;
  wire [4:0] _io_out_T_48_rs2 = _io_out_T_2 == 5'h17 ? io_in[6:2] : _io_out_T_46_rs2;
  wire [4:0] _io_out_T_48_rs3 = _io_out_T_2 == 5'h17 ? io_out_s_0_rs3 : _io_out_T_46_rs3;
  wire [31:0] _io_out_T_50_bits = _io_out_T_2 == 5'h18 ? io_in : _io_out_T_48_bits;
  wire [4:0] _io_out_T_50_rd = _io_out_T_2 == 5'h18 ? io_in[11:7] : _io_out_T_48_rd;
  wire [4:0] _io_out_T_50_rs1 = _io_out_T_2 == 5'h18 ? io_out_s_24_rs1 : _io_out_T_48_rs1;
  wire [4:0] _io_out_T_50_rs2 = _io_out_T_2 == 5'h18 ? io_out_s_24_rs2 : _io_out_T_48_rs2;
  wire [4:0] _io_out_T_50_rs3 = _io_out_T_2 == 5'h18 ? io_out_s_0_rs3 : _io_out_T_48_rs3;
  wire [31:0] _io_out_T_52_bits = _io_out_T_2 == 5'h19 ? io_in : _io_out_T_50_bits;
  wire [4:0] _io_out_T_52_rd = _io_out_T_2 == 5'h19 ? io_in[11:7] : _io_out_T_50_rd;
  wire [4:0] _io_out_T_52_rs1 = _io_out_T_2 == 5'h19 ? io_out_s_24_rs1 : _io_out_T_50_rs1;
  wire [4:0] _io_out_T_52_rs2 = _io_out_T_2 == 5'h19 ? io_out_s_24_rs2 : _io_out_T_50_rs2;
  wire [4:0] _io_out_T_52_rs3 = _io_out_T_2 == 5'h19 ? io_out_s_0_rs3 : _io_out_T_50_rs3;
  wire [31:0] _io_out_T_54_bits = _io_out_T_2 == 5'h1a ? io_in : _io_out_T_52_bits;
  wire [4:0] _io_out_T_54_rd = _io_out_T_2 == 5'h1a ? io_in[11:7] : _io_out_T_52_rd;
  wire [4:0] _io_out_T_54_rs1 = _io_out_T_2 == 5'h1a ? io_out_s_24_rs1 : _io_out_T_52_rs1;
  wire [4:0] _io_out_T_54_rs2 = _io_out_T_2 == 5'h1a ? io_out_s_24_rs2 : _io_out_T_52_rs2;
  wire [4:0] _io_out_T_54_rs3 = _io_out_T_2 == 5'h1a ? io_out_s_0_rs3 : _io_out_T_52_rs3;
  wire [31:0] _io_out_T_56_bits = _io_out_T_2 == 5'h1b ? io_in : _io_out_T_54_bits;
  wire [4:0] _io_out_T_56_rd = _io_out_T_2 == 5'h1b ? io_in[11:7] : _io_out_T_54_rd;
  wire [4:0] _io_out_T_56_rs1 = _io_out_T_2 == 5'h1b ? io_out_s_24_rs1 : _io_out_T_54_rs1;
  wire [4:0] _io_out_T_56_rs2 = _io_out_T_2 == 5'h1b ? io_out_s_24_rs2 : _io_out_T_54_rs2;
  wire [4:0] _io_out_T_56_rs3 = _io_out_T_2 == 5'h1b ? io_out_s_0_rs3 : _io_out_T_54_rs3;
  wire [31:0] _io_out_T_58_bits = _io_out_T_2 == 5'h1c ? io_in : _io_out_T_56_bits;
  wire [4:0] _io_out_T_58_rd = _io_out_T_2 == 5'h1c ? io_in[11:7] : _io_out_T_56_rd;
  wire [4:0] _io_out_T_58_rs1 = _io_out_T_2 == 5'h1c ? io_out_s_24_rs1 : _io_out_T_56_rs1;
  wire [4:0] _io_out_T_58_rs2 = _io_out_T_2 == 5'h1c ? io_out_s_24_rs2 : _io_out_T_56_rs2;
  wire [4:0] _io_out_T_58_rs3 = _io_out_T_2 == 5'h1c ? io_out_s_0_rs3 : _io_out_T_56_rs3;
  wire [31:0] _io_out_T_60_bits = _io_out_T_2 == 5'h1d ? io_in : _io_out_T_58_bits;
  wire [4:0] _io_out_T_60_rd = _io_out_T_2 == 5'h1d ? io_in[11:7] : _io_out_T_58_rd;
  wire [4:0] _io_out_T_60_rs1 = _io_out_T_2 == 5'h1d ? io_out_s_24_rs1 : _io_out_T_58_rs1;
  wire [4:0] _io_out_T_60_rs2 = _io_out_T_2 == 5'h1d ? io_out_s_24_rs2 : _io_out_T_58_rs2;
  wire [4:0] _io_out_T_60_rs3 = _io_out_T_2 == 5'h1d ? io_out_s_0_rs3 : _io_out_T_58_rs3;
  wire [31:0] _io_out_T_62_bits = _io_out_T_2 == 5'h1e ? io_in : _io_out_T_60_bits;
  wire [4:0] _io_out_T_62_rd = _io_out_T_2 == 5'h1e ? io_in[11:7] : _io_out_T_60_rd;
  wire [4:0] _io_out_T_62_rs1 = _io_out_T_2 == 5'h1e ? io_out_s_24_rs1 : _io_out_T_60_rs1;
  wire [4:0] _io_out_T_62_rs2 = _io_out_T_2 == 5'h1e ? io_out_s_24_rs2 : _io_out_T_60_rs2;
  wire [4:0] _io_out_T_62_rs3 = _io_out_T_2 == 5'h1e ? io_out_s_0_rs3 : _io_out_T_60_rs3;
  assign io_out_bits = _io_out_T_2 == 5'h1f ? io_in : _io_out_T_62_bits;
  assign io_out_rd = _io_out_T_2 == 5'h1f ? io_in[11:7] : _io_out_T_62_rd;
  assign io_out_rs1 = _io_out_T_2 == 5'h1f ? io_out_s_24_rs1 : _io_out_T_62_rs1;
  assign io_out_rs2 = _io_out_T_2 == 5'h1f ? io_out_s_24_rs2 : _io_out_T_62_rs2;
  assign io_out_rs3 = _io_out_T_2 == 5'h1f ? io_out_s_0_rs3 : _io_out_T_62_rs3;
  assign io_rvc = io_in[1:0] != 2'h3;
endmodule